/*
 * Copyright (c) 2018 Sprocket
 *
 * This is free software: you can redistribute it and/or modify
 * it under the terms of the GNU Affero General Public License with
 * additional permissions to the one published by the Free Software
 * Foundation, either version 3 of the License, or (at your option)
 * any later version. For more information see LICENSE.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU Affero General Public License for more details.
 *
 * You should have received a copy of the GNU Affero General Public License
 * along with this program. If not, see <http://www.gnu.org/licenses/>.
 */

module JH512 (
	input clk,
	input [1023:0] state,
	input [127:0] data,
	output [511:0] hash
);

	reg [127:0] data_le;

	reg [127:0] d00,d01,d02,d03,d04,d05,d06,d07,d08,d09;
	reg [127:0] d10,d11,d12,d13,d14,d15,d16,d17,d18,d19;
	reg [127:0] d20,d21,d22,d23,d24,d25,d26,d27,d28,d29;
	reg [127:0] d30,d31,d32,d33,d34,d35,d36,d37,d38,d39;
	reg [127:0] d40,d41,d42,d43,d44,d45;

	reg [1023:0] H00, H01, H10, H11;
	reg [511:0]  H20, H21;
	assign hash = H21;
	
	wire [1023:0] state0, state1;
	
	F8 F8_0 (clk, H01, state0);
	F8 F8_1 (clk, H11, state1);

	always @ ( posedge clk ) begin

		data_le <= { // 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080,
						data[  7:  0],
						data[ 15:  8],
						data[ 23: 16],
						data[ 31: 24],
						data[ 39: 32],
						data[ 47: 40],
						data[ 55: 48],
						data[ 63: 56],
						data[ 71: 64],
						data[ 79: 72],
						data[ 87: 80],
						data[ 95: 88],
						data[103: 96],
						data[111:104],
						data[119:112],
						data[127:120] };

		H00 <= state;

		H01[1023:136] <= H00[1023:136];
		H01[ 135:128] <= H00[ 135:128] ^ 8'h80;
		H01[ 127:  0] <= H00[ 127:  0] ^ data_le[127:0];

		H10 <= state0;

		H11[1023:648] <= H10[1023:648];
		H11[ 647:640] <= H10[ 647:640] ^ 8'h80;
		H11[ 639:512] <= H10[ 639:512] ^ d45;
		H11[ 511:496] <= H10[ 511:496] ^ 16'h8002;
		H11[ 495:  0] <= H10[ 495:  0];

//		data1 <= 512'h80020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

		H20 <= state1[1023:512];

		H21[  7:  0] <= H20[511:504] ^ 8'h80;
		H21[ 15:  8] <= H20[503:496] ^ 8'h02;
		H21[ 23: 16] <= H20[495:488];
		H21[ 31: 24] <= H20[487:480];
		H21[ 39: 32] <= H20[479:472];
		H21[ 47: 40] <= H20[471:464];
		H21[ 55: 48] <= H20[463:456];
		H21[ 63: 56] <= H20[455:448];
		H21[ 71: 64] <= H20[447:440];
		H21[ 79: 72] <= H20[439:432];
		H21[ 87: 80] <= H20[431:424];
		H21[ 95: 88] <= H20[423:416];
		H21[103: 96] <= H20[415:408];
		H21[111:104] <= H20[407:400];
		H21[119:112] <= H20[399:392];
		H21[127:120] <= H20[391:384];
		H21[135:128] <= H20[383:376];
		H21[143:136] <= H20[375:368];
		H21[151:144] <= H20[367:360];
		H21[159:152] <= H20[359:352];
		H21[167:160] <= H20[351:344];
		H21[175:168] <= H20[343:336];
		H21[183:176] <= H20[335:328];
		H21[191:184] <= H20[327:320];
		H21[199:192] <= H20[319:312];
		H21[207:200] <= H20[311:304];
		H21[215:208] <= H20[303:296];
		H21[223:216] <= H20[295:288];
		H21[231:224] <= H20[287:280];
		H21[239:232] <= H20[279:272];
		H21[247:240] <= H20[271:264];
		H21[255:248] <= H20[263:256];
		H21[263:256] <= H20[255:248];
		H21[271:264] <= H20[247:240];
		H21[279:272] <= H20[239:232];
		H21[287:280] <= H20[231:224];
		H21[295:288] <= H20[223:216];
		H21[303:296] <= H20[215:208];
		H21[311:304] <= H20[207:200];
		H21[319:312] <= H20[199:192];
		H21[327:320] <= H20[191:184];
		H21[335:328] <= H20[183:176];
		H21[343:336] <= H20[175:168];
		H21[351:344] <= H20[167:160];
		H21[359:352] <= H20[159:152];
		H21[367:360] <= H20[151:144];
		H21[375:368] <= H20[143:136];
		H21[383:376] <= H20[135:128];
		H21[391:384] <= H20[127:120];
		H21[399:392] <= H20[119:112];
		H21[407:400] <= H20[111:104];
		H21[415:408] <= H20[103: 96];
		H21[423:416] <= H20[ 95: 88];
		H21[431:424] <= H20[ 87: 80];
		H21[439:432] <= H20[ 79: 72];
		H21[447:440] <= H20[ 71: 64];
		H21[455:448] <= H20[ 63: 56];
		H21[463:456] <= H20[ 55: 48];
		H21[471:464] <= H20[ 47: 40];
		H21[479:472] <= H20[ 39: 32];
		H21[487:480] <= H20[ 31: 24];
		H21[495:488] <= H20[ 23: 16];
		H21[503:496] <= H20[ 15:  8];
		H21[511:504] <= H20[  7:  0];

		d45 <= d44;
		d44 <= d43;
		d43 <= d42;
		d42 <= d41;
		d41 <= d40;
		d40 <= d39;
		d39 <= d38;
		d38 <= d37;
		d37 <= d36;
		d36 <= d35;
		d35 <= d34;
		d34 <= d33;
		d33 <= d32;
		d32 <= d31;
		d31 <= d30;
		d30 <= d29;
		d29 <= d28;
		d28 <= d27;
		d27 <= d26;
		d26 <= d25;
		d25 <= d24;
		d24 <= d23;
		d23 <= d22;
		d22 <= d21;
		d21 <= d20;
		d20 <= d19;
		d19 <= d18;
		d18 <= d17;
		d17 <= d16;
		d16 <= d15;
		d15 <= d14;
		d14 <= d13;
		d13 <= d12;
		d12 <= d11;
		d11 <= d10;
		d10 <= d09;
		d09 <= d08;
		d08 <= d07;
		d07 <= d06;
		d06 <= d05;
		d05 <= d04;
		d04 <= d03;
		d03 <= d02;
		d02 <= d01;
		d01 <= d00;
		d00 <= data_le[127:0];

	end
	
endmodule

module F8 (
	input clk,
	input [1023:0] state_in,
	output reg [1023:0] state_out
);

	reg [255:0] R;
	reg [1023:0] i;
	wire [1023:0] i0,f0;

	wire [1023:0] a00,a01,a02,a03,a04,a05,a06,a07,a08,a09;
	wire [1023:0] a10,a11,a12,a13,a14,a15,a16,a17,a18,a19;
	wire [1023:0] a20,a21,a22,a23,a24,a25,a26,a27,a28,a29;
	wire [1023:0] a30,a31,a32,a33,a34,a35,a36,a37,a38,a39,a40,a41;
	
	wire [255:0] r00,r01,r02,r03,r04,r05,r06,r07,r08,r09;
	wire [255:0] r10,r11,r12,r13,r14,r15,r16,r17,r18,r19;
	wire [255:0] r20,r21,r22,r23,r24,r25,r26,r27,r28,r29;
	wire [255:0] r30,r31,r32,r33,r34,r35,r36,r37,r38,r39,r40,r41;

	reg [1023:0] a00x,a01x,a02x,a03x,a04x,a05x,a06x,a07x,a08x,a09x;
	reg [1023:0] a10x,a11x,a12x,a13x,a14x,a15x,a16x,a17x,a18x,a19x;
	reg [1023:0] a20x,a21x,a22x,a23x,a24x,a25x,a26x,a27x,a28x,a29x;
	reg [1023:0] a30x,a31x,a32x,a33x,a34x,a35x,a36x,a37x,a38x,a39x,a40x,a41x;
	
	reg [255:0] r00x,r01x,r02x,r03x,r04x,r05x,r06x,r07x,r08x,r09x;
	reg [255:0] r10x,r11x,r12x,r13x,r14x,r15x,r16x,r17x,r18x,r19x;
	reg [255:0] r20x,r21x,r22x,r23x,r24x,r25x,r26x,r27x,r28x,r29x;
	reg [255:0] r30x,r31x,r32x,r33x,r34x,r35x,r36x,r37x,r38x,r39x,r40x,r41x;
	
	jh_init jh_init  (i,i0);
	jh_round_a jh00a (i0, R, a00);
	jh_round_b jh00b (    R, r00);
	jh_round_a jh01a (a00x,r00x,a01);
	jh_round_b jh01b (    r00x,r01);
	jh_round_a jh02a (a01x,r01x,a02);
	jh_round_b jh02b (    r01x,r02);
	jh_round_a jh03a (a02x,r02x,a03);
	jh_round_b jh03b (    r02x,r03);
	jh_round_a jh04a (a03x,r03x,a04);
	jh_round_b jh04b (    r03x,r04);
	jh_round_a jh05a (a04x,r04x,a05);
	jh_round_b jh05b (    r04x,r05);
	jh_round_a jh06a (a05x,r05x,a06);
	jh_round_b jh06b (    r05x,r06);
	jh_round_a jh07a (a06x,r06x,a07);
	jh_round_b jh07b (    r06x,r07);
	jh_round_a jh08a (a07x,r07x,a08);
	jh_round_b jh08b (    r07x,r08);
	jh_round_a jh09a (a08x,r08x,a09);
	jh_round_b jh09b (    r08x,r09);
	jh_round_a jh10a (a09x,r09x,a10);
	jh_round_b jh10b (    r09x,r10);
	jh_round_a jh11a (a10x,r10x,a11);
	jh_round_b jh11b (    r10x,r11);
	jh_round_a jh12a (a11x,r11x,a12);
	jh_round_b jh12b (    r11x,r12);
	jh_round_a jh13a (a12x,r12x,a13);
	jh_round_b jh13b (    r12x,r13);
	jh_round_a jh14a (a13x,r13x,a14);
	jh_round_b jh14b (    r13x,r14);
	jh_round_a jh15a (a14x,r14x,a15);
	jh_round_b jh15b (    r14x,r15);
	jh_round_a jh16a (a15x,r15x,a16);
	jh_round_b jh16b (    r15x,r16);
	jh_round_a jh17a (a16x,r16x,a17);
	jh_round_b jh17b (    r16x,r17);
	jh_round_a jh18a (a17x,r17x,a18);
	jh_round_b jh18b (    r17x,r18);
	jh_round_a jh19a (a18x,r18x,a19);
	jh_round_b jh19b (    r18x,r19);
	jh_round_a jh20a (a19x,r19x,a20);
	jh_round_b jh20b (    r19x,r20);
	jh_round_a jh21a (a20x,r20x,a21);
	jh_round_b jh21b (    r20x,r21);
	jh_round_a jh22a (a21x,r21x,a22);
	jh_round_b jh22b (    r21x,r22);
	jh_round_a jh23a (a22x,r22x,a23);
	jh_round_b jh23b (    r22x,r23);
	jh_round_a jh24a (a23x,r23x,a24);
	jh_round_b jh24b (    r23x,r24);
	jh_round_a jh25a (a24x,r24x,a25);
	jh_round_b jh25b (    r24x,r25);
	jh_round_a jh26a (a25x,r25x,a26);
	jh_round_b jh26b (    r25x,r26);
	jh_round_a jh27a (a26x,r26x,a27);
	jh_round_b jh27b (    r26x,r27);
	jh_round_a jh28a (a27x,r27x,a28);
	jh_round_b jh28b (    r27x,r28);
	jh_round_a jh29a (a28x,r28x,a29);
	jh_round_b jh29b (    r28x,r29);
	jh_round_a jh30a (a29x,r29x,a30);
	jh_round_b jh30b (    r29x,r30);
	jh_round_a jh31a (a30x,r30x,a31);
	jh_round_b jh31b (    r30x,r31);
	jh_round_a jh32a (a31x,r31x,a32);
	jh_round_b jh32b (    r31x,r32);
	jh_round_a jh33a (a32x,r32x,a33);
	jh_round_b jh33b (    r32x,r33);
	jh_round_a jh34a (a33x,r33x,a34);
	jh_round_b jh34b (    r33x,r34);
	jh_round_a jh35a (a34x,r34x,a35);
	jh_round_b jh35b (    r34x,r35);
	jh_round_a jh36a (a35x,r35x,a36);
	jh_round_b jh36b (    r35x,r36);
	jh_round_a jh37a (a36x,r36x,a37);
	jh_round_b jh37b (    r36x,r37);
	jh_round_a jh38a (a37x,r37x,a38);
	jh_round_b jh38b (    r37x,r38);
	jh_round_a jh39a (a38x,r38x,a39);
	jh_round_b jh39b (    r38x,r39);
	jh_round_a jh40a (a39x,r39x,a40);
	jh_round_b jh40b (    r39x,r40);
	jh_round_a jh41a (a40x,r40x,a41);
//	jh_round_b jh41b (    r40,r41);
	jh_final jh_final(a41x,f0);

	always @ ( posedge clk ) begin
	
		i <= state_in;
		R <= 256'h544ce660d09af45b990aee48ae837b5c7cbea95766c8df4d10933dcfe6679056;
		state_out <= f0;
		
		a00x <= a00;
		r00x <= r00;
		a01x <= a01;
		r01x <= r01;
		a02x <= a02;
		r02x <= r02;
		a03x <= a03;
		r03x <= r03;
		a04x <= a04;
		r04x <= r04;
		a05x <= a05;
		r05x <= r05;
		a06x <= a06;
		r06x <= r06;
		a07x <= a07;
		r07x <= r07;
		a08x <= a08;
		r08x <= r08;
		a09x <= a09;
		r09x <= r09;
		a10x <= a10;
		r10x <= r10;
		a11x <= a11;
		r11x <= r11;
		a12x <= a12;
		r12x <= r12;
		a13x <= a13;
		r13x <= r13;
		a14x <= a14;
		r14x <= r14;
		a15x <= a15;
		r15x <= r15;
		a16x <= a16;
		r16x <= r16;
		a17x <= a17;
		r17x <= r17;
		a18x <= a18;
		r18x <= r18;
		a19x <= a19;
		r19x <= r19;
		a20x <= a20;
		r20x <= r20;
		a21x <= a21;
		r21x <= r21;
		a22x <= a22;
		r22x <= r22;
		a23x <= a23;
		r23x <= r23;
		a24x <= a24;
		r24x <= r24;
		a25x <= a25;
		r25x <= r25;
		a26x <= a26;
		r26x <= r26;
		a27x <= a27;
		r27x <= r27;
		a28x <= a28;
		r28x <= r28;
		a29x <= a29;
		r29x <= r29;
		a30x <= a30;
		r30x <= r30;
		a31x <= a31;
		r31x <= r31;
		a32x <= a32;
		r32x <= r32;
		a33x <= a33;
		r33x <= r33;
		a34x <= a34;
		r34x <= r34;
		a35x <= a35;
		r35x <= r35;
		a36x <= a36;
		r36x <= r36;
		a37x <= a37;
		r37x <= r37;
		a38x <= a38;
		r38x <= r38;
		a39x <= a39;
		r39x <= r39;
		a40x <= a40;
		r40x <= r40;
		a41x <= a41;
		r41x <= r41;

	end
	
endmodule


module jh_init (
	input [1023:0] in,
	output [1023:0] out
);

	assign out[3:0] = { in[7], in[263], in[519], in[775] };
	assign out[11:8] = { in[6], in[262], in[518], in[774] };
	assign out[19:16] = { in[5], in[261], in[517], in[773] };
	assign out[27:24] = { in[4], in[260], in[516], in[772] };
	assign out[35:32] = { in[3], in[259], in[515], in[771] };
	assign out[43:40] = { in[2], in[258], in[514], in[770] };
	assign out[51:48] = { in[1], in[257], in[513], in[769] };
	assign out[59:56] = { in[0], in[256], in[512], in[768] };
	assign out[67:64] = { in[15], in[271], in[527], in[783] };
	assign out[75:72] = { in[14], in[270], in[526], in[782] };
	assign out[83:80] = { in[13], in[269], in[525], in[781] };
	assign out[91:88] = { in[12], in[268], in[524], in[780] };
	assign out[99:96] = { in[11], in[267], in[523], in[779] };
	assign out[107:104] = { in[10], in[266], in[522], in[778] };
	assign out[115:112] = { in[9], in[265], in[521], in[777] };
	assign out[123:120] = { in[8], in[264], in[520], in[776] };
	assign out[131:128] = { in[23], in[279], in[535], in[791] };
	assign out[139:136] = { in[22], in[278], in[534], in[790] };
	assign out[147:144] = { in[21], in[277], in[533], in[789] };
	assign out[155:152] = { in[20], in[276], in[532], in[788] };
	assign out[163:160] = { in[19], in[275], in[531], in[787] };
	assign out[171:168] = { in[18], in[274], in[530], in[786] };
	assign out[179:176] = { in[17], in[273], in[529], in[785] };
	assign out[187:184] = { in[16], in[272], in[528], in[784] };
	assign out[195:192] = { in[31], in[287], in[543], in[799] };
	assign out[203:200] = { in[30], in[286], in[542], in[798] };
	assign out[211:208] = { in[29], in[285], in[541], in[797] };
	assign out[219:216] = { in[28], in[284], in[540], in[796] };
	assign out[227:224] = { in[27], in[283], in[539], in[795] };
	assign out[235:232] = { in[26], in[282], in[538], in[794] };
	assign out[243:240] = { in[25], in[281], in[537], in[793] };
	assign out[251:248] = { in[24], in[280], in[536], in[792] };
	assign out[259:256] = { in[39], in[295], in[551], in[807] };
	assign out[267:264] = { in[38], in[294], in[550], in[806] };
	assign out[275:272] = { in[37], in[293], in[549], in[805] };
	assign out[283:280] = { in[36], in[292], in[548], in[804] };
	assign out[291:288] = { in[35], in[291], in[547], in[803] };
	assign out[299:296] = { in[34], in[290], in[546], in[802] };
	assign out[307:304] = { in[33], in[289], in[545], in[801] };
	assign out[315:312] = { in[32], in[288], in[544], in[800] };
	assign out[323:320] = { in[47], in[303], in[559], in[815] };
	assign out[331:328] = { in[46], in[302], in[558], in[814] };
	assign out[339:336] = { in[45], in[301], in[557], in[813] };
	assign out[347:344] = { in[44], in[300], in[556], in[812] };
	assign out[355:352] = { in[43], in[299], in[555], in[811] };
	assign out[363:360] = { in[42], in[298], in[554], in[810] };
	assign out[371:368] = { in[41], in[297], in[553], in[809] };
	assign out[379:376] = { in[40], in[296], in[552], in[808] };
	assign out[387:384] = { in[55], in[311], in[567], in[823] };
	assign out[395:392] = { in[54], in[310], in[566], in[822] };
	assign out[403:400] = { in[53], in[309], in[565], in[821] };
	assign out[411:408] = { in[52], in[308], in[564], in[820] };
	assign out[419:416] = { in[51], in[307], in[563], in[819] };
	assign out[427:424] = { in[50], in[306], in[562], in[818] };
	assign out[435:432] = { in[49], in[305], in[561], in[817] };
	assign out[443:440] = { in[48], in[304], in[560], in[816] };
	assign out[451:448] = { in[63], in[319], in[575], in[831] };
	assign out[459:456] = { in[62], in[318], in[574], in[830] };
	assign out[467:464] = { in[61], in[317], in[573], in[829] };
	assign out[475:472] = { in[60], in[316], in[572], in[828] };
	assign out[483:480] = { in[59], in[315], in[571], in[827] };
	assign out[491:488] = { in[58], in[314], in[570], in[826] };
	assign out[499:496] = { in[57], in[313], in[569], in[825] };
	assign out[507:504] = { in[56], in[312], in[568], in[824] };
	assign out[515:512] = { in[71], in[327], in[583], in[839] };
	assign out[523:520] = { in[70], in[326], in[582], in[838] };
	assign out[531:528] = { in[69], in[325], in[581], in[837] };
	assign out[539:536] = { in[68], in[324], in[580], in[836] };
	assign out[547:544] = { in[67], in[323], in[579], in[835] };
	assign out[555:552] = { in[66], in[322], in[578], in[834] };
	assign out[563:560] = { in[65], in[321], in[577], in[833] };
	assign out[571:568] = { in[64], in[320], in[576], in[832] };
	assign out[579:576] = { in[79], in[335], in[591], in[847] };
	assign out[587:584] = { in[78], in[334], in[590], in[846] };
	assign out[595:592] = { in[77], in[333], in[589], in[845] };
	assign out[603:600] = { in[76], in[332], in[588], in[844] };
	assign out[611:608] = { in[75], in[331], in[587], in[843] };
	assign out[619:616] = { in[74], in[330], in[586], in[842] };
	assign out[627:624] = { in[73], in[329], in[585], in[841] };
	assign out[635:632] = { in[72], in[328], in[584], in[840] };
	assign out[643:640] = { in[87], in[343], in[599], in[855] };
	assign out[651:648] = { in[86], in[342], in[598], in[854] };
	assign out[659:656] = { in[85], in[341], in[597], in[853] };
	assign out[667:664] = { in[84], in[340], in[596], in[852] };
	assign out[675:672] = { in[83], in[339], in[595], in[851] };
	assign out[683:680] = { in[82], in[338], in[594], in[850] };
	assign out[691:688] = { in[81], in[337], in[593], in[849] };
	assign out[699:696] = { in[80], in[336], in[592], in[848] };
	assign out[707:704] = { in[95], in[351], in[607], in[863] };
	assign out[715:712] = { in[94], in[350], in[606], in[862] };
	assign out[723:720] = { in[93], in[349], in[605], in[861] };
	assign out[731:728] = { in[92], in[348], in[604], in[860] };
	assign out[739:736] = { in[91], in[347], in[603], in[859] };
	assign out[747:744] = { in[90], in[346], in[602], in[858] };
	assign out[755:752] = { in[89], in[345], in[601], in[857] };
	assign out[763:760] = { in[88], in[344], in[600], in[856] };
	assign out[771:768] = { in[103], in[359], in[615], in[871] };
	assign out[779:776] = { in[102], in[358], in[614], in[870] };
	assign out[787:784] = { in[101], in[357], in[613], in[869] };
	assign out[795:792] = { in[100], in[356], in[612], in[868] };
	assign out[803:800] = { in[99], in[355], in[611], in[867] };
	assign out[811:808] = { in[98], in[354], in[610], in[866] };
	assign out[819:816] = { in[97], in[353], in[609], in[865] };
	assign out[827:824] = { in[96], in[352], in[608], in[864] };
	assign out[835:832] = { in[111], in[367], in[623], in[879] };
	assign out[843:840] = { in[110], in[366], in[622], in[878] };
	assign out[851:848] = { in[109], in[365], in[621], in[877] };
	assign out[859:856] = { in[108], in[364], in[620], in[876] };
	assign out[867:864] = { in[107], in[363], in[619], in[875] };
	assign out[875:872] = { in[106], in[362], in[618], in[874] };
	assign out[883:880] = { in[105], in[361], in[617], in[873] };
	assign out[891:888] = { in[104], in[360], in[616], in[872] };
	assign out[899:896] = { in[119], in[375], in[631], in[887] };
	assign out[907:904] = { in[118], in[374], in[630], in[886] };
	assign out[915:912] = { in[117], in[373], in[629], in[885] };
	assign out[923:920] = { in[116], in[372], in[628], in[884] };
	assign out[931:928] = { in[115], in[371], in[627], in[883] };
	assign out[939:936] = { in[114], in[370], in[626], in[882] };
	assign out[947:944] = { in[113], in[369], in[625], in[881] };
	assign out[955:952] = { in[112], in[368], in[624], in[880] };
	assign out[963:960] = { in[127], in[383], in[639], in[895] };
	assign out[971:968] = { in[126], in[382], in[638], in[894] };
	assign out[979:976] = { in[125], in[381], in[637], in[893] };
	assign out[987:984] = { in[124], in[380], in[636], in[892] };
	assign out[995:992] = { in[123], in[379], in[635], in[891] };
	assign out[1003:1000] = { in[122], in[378], in[634], in[890] };
	assign out[1011:1008] = { in[121], in[377], in[633], in[889] };
	assign out[1019:1016] = { in[120], in[376], in[632], in[888] };
	assign out[7:4] = { in[135], in[391], in[647], in[903] };
	assign out[15:12] = { in[134], in[390], in[646], in[902] };
	assign out[23:20] = { in[133], in[389], in[645], in[901] };
	assign out[31:28] = { in[132], in[388], in[644], in[900] };
	assign out[39:36] = { in[131], in[387], in[643], in[899] };
	assign out[47:44] = { in[130], in[386], in[642], in[898] };
	assign out[55:52] = { in[129], in[385], in[641], in[897] };
	assign out[63:60] = { in[128], in[384], in[640], in[896] };
	assign out[71:68] = { in[143], in[399], in[655], in[911] };
	assign out[79:76] = { in[142], in[398], in[654], in[910] };
	assign out[87:84] = { in[141], in[397], in[653], in[909] };
	assign out[95:92] = { in[140], in[396], in[652], in[908] };
	assign out[103:100] = { in[139], in[395], in[651], in[907] };
	assign out[111:108] = { in[138], in[394], in[650], in[906] };
	assign out[119:116] = { in[137], in[393], in[649], in[905] };
	assign out[127:124] = { in[136], in[392], in[648], in[904] };
	assign out[135:132] = { in[151], in[407], in[663], in[919] };
	assign out[143:140] = { in[150], in[406], in[662], in[918] };
	assign out[151:148] = { in[149], in[405], in[661], in[917] };
	assign out[159:156] = { in[148], in[404], in[660], in[916] };
	assign out[167:164] = { in[147], in[403], in[659], in[915] };
	assign out[175:172] = { in[146], in[402], in[658], in[914] };
	assign out[183:180] = { in[145], in[401], in[657], in[913] };
	assign out[191:188] = { in[144], in[400], in[656], in[912] };
	assign out[199:196] = { in[159], in[415], in[671], in[927] };
	assign out[207:204] = { in[158], in[414], in[670], in[926] };
	assign out[215:212] = { in[157], in[413], in[669], in[925] };
	assign out[223:220] = { in[156], in[412], in[668], in[924] };
	assign out[231:228] = { in[155], in[411], in[667], in[923] };
	assign out[239:236] = { in[154], in[410], in[666], in[922] };
	assign out[247:244] = { in[153], in[409], in[665], in[921] };
	assign out[255:252] = { in[152], in[408], in[664], in[920] };
	assign out[263:260] = { in[167], in[423], in[679], in[935] };
	assign out[271:268] = { in[166], in[422], in[678], in[934] };
	assign out[279:276] = { in[165], in[421], in[677], in[933] };
	assign out[287:284] = { in[164], in[420], in[676], in[932] };
	assign out[295:292] = { in[163], in[419], in[675], in[931] };
	assign out[303:300] = { in[162], in[418], in[674], in[930] };
	assign out[311:308] = { in[161], in[417], in[673], in[929] };
	assign out[319:316] = { in[160], in[416], in[672], in[928] };
	assign out[327:324] = { in[175], in[431], in[687], in[943] };
	assign out[335:332] = { in[174], in[430], in[686], in[942] };
	assign out[343:340] = { in[173], in[429], in[685], in[941] };
	assign out[351:348] = { in[172], in[428], in[684], in[940] };
	assign out[359:356] = { in[171], in[427], in[683], in[939] };
	assign out[367:364] = { in[170], in[426], in[682], in[938] };
	assign out[375:372] = { in[169], in[425], in[681], in[937] };
	assign out[383:380] = { in[168], in[424], in[680], in[936] };
	assign out[391:388] = { in[183], in[439], in[695], in[951] };
	assign out[399:396] = { in[182], in[438], in[694], in[950] };
	assign out[407:404] = { in[181], in[437], in[693], in[949] };
	assign out[415:412] = { in[180], in[436], in[692], in[948] };
	assign out[423:420] = { in[179], in[435], in[691], in[947] };
	assign out[431:428] = { in[178], in[434], in[690], in[946] };
	assign out[439:436] = { in[177], in[433], in[689], in[945] };
	assign out[447:444] = { in[176], in[432], in[688], in[944] };
	assign out[455:452] = { in[191], in[447], in[703], in[959] };
	assign out[463:460] = { in[190], in[446], in[702], in[958] };
	assign out[471:468] = { in[189], in[445], in[701], in[957] };
	assign out[479:476] = { in[188], in[444], in[700], in[956] };
	assign out[487:484] = { in[187], in[443], in[699], in[955] };
	assign out[495:492] = { in[186], in[442], in[698], in[954] };
	assign out[503:500] = { in[185], in[441], in[697], in[953] };
	assign out[511:508] = { in[184], in[440], in[696], in[952] };
	assign out[519:516] = { in[199], in[455], in[711], in[967] };
	assign out[527:524] = { in[198], in[454], in[710], in[966] };
	assign out[535:532] = { in[197], in[453], in[709], in[965] };
	assign out[543:540] = { in[196], in[452], in[708], in[964] };
	assign out[551:548] = { in[195], in[451], in[707], in[963] };
	assign out[559:556] = { in[194], in[450], in[706], in[962] };
	assign out[567:564] = { in[193], in[449], in[705], in[961] };
	assign out[575:572] = { in[192], in[448], in[704], in[960] };
	assign out[583:580] = { in[207], in[463], in[719], in[975] };
	assign out[591:588] = { in[206], in[462], in[718], in[974] };
	assign out[599:596] = { in[205], in[461], in[717], in[973] };
	assign out[607:604] = { in[204], in[460], in[716], in[972] };
	assign out[615:612] = { in[203], in[459], in[715], in[971] };
	assign out[623:620] = { in[202], in[458], in[714], in[970] };
	assign out[631:628] = { in[201], in[457], in[713], in[969] };
	assign out[639:636] = { in[200], in[456], in[712], in[968] };
	assign out[647:644] = { in[215], in[471], in[727], in[983] };
	assign out[655:652] = { in[214], in[470], in[726], in[982] };
	assign out[663:660] = { in[213], in[469], in[725], in[981] };
	assign out[671:668] = { in[212], in[468], in[724], in[980] };
	assign out[679:676] = { in[211], in[467], in[723], in[979] };
	assign out[687:684] = { in[210], in[466], in[722], in[978] };
	assign out[695:692] = { in[209], in[465], in[721], in[977] };
	assign out[703:700] = { in[208], in[464], in[720], in[976] };
	assign out[711:708] = { in[223], in[479], in[735], in[991] };
	assign out[719:716] = { in[222], in[478], in[734], in[990] };
	assign out[727:724] = { in[221], in[477], in[733], in[989] };
	assign out[735:732] = { in[220], in[476], in[732], in[988] };
	assign out[743:740] = { in[219], in[475], in[731], in[987] };
	assign out[751:748] = { in[218], in[474], in[730], in[986] };
	assign out[759:756] = { in[217], in[473], in[729], in[985] };
	assign out[767:764] = { in[216], in[472], in[728], in[984] };
	assign out[775:772] = { in[231], in[487], in[743], in[999] };
	assign out[783:780] = { in[230], in[486], in[742], in[998] };
	assign out[791:788] = { in[229], in[485], in[741], in[997] };
	assign out[799:796] = { in[228], in[484], in[740], in[996] };
	assign out[807:804] = { in[227], in[483], in[739], in[995] };
	assign out[815:812] = { in[226], in[482], in[738], in[994] };
	assign out[823:820] = { in[225], in[481], in[737], in[993] };
	assign out[831:828] = { in[224], in[480], in[736], in[992] };
	assign out[839:836] = { in[239], in[495], in[751], in[1007] };
	assign out[847:844] = { in[238], in[494], in[750], in[1006] };
	assign out[855:852] = { in[237], in[493], in[749], in[1005] };
	assign out[863:860] = { in[236], in[492], in[748], in[1004] };
	assign out[871:868] = { in[235], in[491], in[747], in[1003] };
	assign out[879:876] = { in[234], in[490], in[746], in[1002] };
	assign out[887:884] = { in[233], in[489], in[745], in[1001] };
	assign out[895:892] = { in[232], in[488], in[744], in[1000] };
	assign out[903:900] = { in[247], in[503], in[759], in[1015] };
	assign out[911:908] = { in[246], in[502], in[758], in[1014] };
	assign out[919:916] = { in[245], in[501], in[757], in[1013] };
	assign out[927:924] = { in[244], in[500], in[756], in[1012] };
	assign out[935:932] = { in[243], in[499], in[755], in[1011] };
	assign out[943:940] = { in[242], in[498], in[754], in[1010] };
	assign out[951:948] = { in[241], in[497], in[753], in[1009] };
	assign out[959:956] = { in[240], in[496], in[752], in[1008] };
	assign out[967:964] = { in[255], in[511], in[767], in[1023] };
	assign out[975:972] = { in[254], in[510], in[766], in[1022] };
	assign out[983:980] = { in[253], in[509], in[765], in[1021] };
	assign out[991:988] = { in[252], in[508], in[764], in[1020] };
	assign out[999:996] = { in[251], in[507], in[763], in[1019] };
	assign out[1007:1004] = { in[250], in[506], in[762], in[1018] };
	assign out[1015:1012] = { in[249], in[505], in[761], in[1017] };
	assign out[1023:1020] = { in[248], in[504], in[760], in[1016] };
	
endmodule

module jh_round_a (
	input [1023:0] state_in,
	input [255:0] round_in,
	output [1023:0] out
);         

	wire [3:0] sbox [0:31] = { 4'h9,4'h0,4'h4,4'hb,4'hd,4'hc,4'h3,4'hf,4'h1,4'ha,4'h2,4'h6,4'h7,4'h5,4'h8,4'he,4'h3,4'hc,4'h6,4'hd,4'h5,4'h7,4'h1,4'h9,4'hf,4'h2,4'h0,4'h4,4'hb,4'ha,4'he,4'h8 };
	
	wire [1023:0] L1;

	assign L1[1023:1020] = sbox[ { round_in[255], state_in[1023:1020] } ];
	assign L1[1019:1016] = sbox[ { round_in[254], state_in[1019:1016] } ];
	assign L1[1015:1012] = sbox[ { round_in[253], state_in[1015:1012] } ];
	assign L1[1011:1008] = sbox[ { round_in[252], state_in[1011:1008] } ];
	assign L1[1007:1004] = sbox[ { round_in[251], state_in[1007:1004] } ];
	assign L1[1003:1000] = sbox[ { round_in[250], state_in[1003:1000] } ];
	assign L1[999:996] = sbox[ { round_in[249], state_in[999:996] } ];
	assign L1[995:992] = sbox[ { round_in[248], state_in[995:992] } ];
	assign L1[991:988] = sbox[ { round_in[247], state_in[991:988] } ];
	assign L1[987:984] = sbox[ { round_in[246], state_in[987:984] } ];
	assign L1[983:980] = sbox[ { round_in[245], state_in[983:980] } ];
	assign L1[979:976] = sbox[ { round_in[244], state_in[979:976] } ];
	assign L1[975:972] = sbox[ { round_in[243], state_in[975:972] } ];
	assign L1[971:968] = sbox[ { round_in[242], state_in[971:968] } ];
	assign L1[967:964] = sbox[ { round_in[241], state_in[967:964] } ];
	assign L1[963:960] = sbox[ { round_in[240], state_in[963:960] } ];
	assign L1[959:956] = sbox[ { round_in[239], state_in[959:956] } ];
	assign L1[955:952] = sbox[ { round_in[238], state_in[955:952] } ];
	assign L1[951:948] = sbox[ { round_in[237], state_in[951:948] } ];
	assign L1[947:944] = sbox[ { round_in[236], state_in[947:944] } ];
	assign L1[943:940] = sbox[ { round_in[235], state_in[943:940] } ];
	assign L1[939:936] = sbox[ { round_in[234], state_in[939:936] } ];
	assign L1[935:932] = sbox[ { round_in[233], state_in[935:932] } ];
	assign L1[931:928] = sbox[ { round_in[232], state_in[931:928] } ];
	assign L1[927:924] = sbox[ { round_in[231], state_in[927:924] } ];
	assign L1[923:920] = sbox[ { round_in[230], state_in[923:920] } ];
	assign L1[919:916] = sbox[ { round_in[229], state_in[919:916] } ];
	assign L1[915:912] = sbox[ { round_in[228], state_in[915:912] } ];
	assign L1[911:908] = sbox[ { round_in[227], state_in[911:908] } ];
	assign L1[907:904] = sbox[ { round_in[226], state_in[907:904] } ];
	assign L1[903:900] = sbox[ { round_in[225], state_in[903:900] } ];
	assign L1[899:896] = sbox[ { round_in[224], state_in[899:896] } ];
	assign L1[895:892] = sbox[ { round_in[223], state_in[895:892] } ];
	assign L1[891:888] = sbox[ { round_in[222], state_in[891:888] } ];
	assign L1[887:884] = sbox[ { round_in[221], state_in[887:884] } ];
	assign L1[883:880] = sbox[ { round_in[220], state_in[883:880] } ];
	assign L1[879:876] = sbox[ { round_in[219], state_in[879:876] } ];
	assign L1[875:872] = sbox[ { round_in[218], state_in[875:872] } ];
	assign L1[871:868] = sbox[ { round_in[217], state_in[871:868] } ];
	assign L1[867:864] = sbox[ { round_in[216], state_in[867:864] } ];
	assign L1[863:860] = sbox[ { round_in[215], state_in[863:860] } ];
	assign L1[859:856] = sbox[ { round_in[214], state_in[859:856] } ];
	assign L1[855:852] = sbox[ { round_in[213], state_in[855:852] } ];
	assign L1[851:848] = sbox[ { round_in[212], state_in[851:848] } ];
	assign L1[847:844] = sbox[ { round_in[211], state_in[847:844] } ];
	assign L1[843:840] = sbox[ { round_in[210], state_in[843:840] } ];
	assign L1[839:836] = sbox[ { round_in[209], state_in[839:836] } ];
	assign L1[835:832] = sbox[ { round_in[208], state_in[835:832] } ];
	assign L1[831:828] = sbox[ { round_in[207], state_in[831:828] } ];
	assign L1[827:824] = sbox[ { round_in[206], state_in[827:824] } ];
	assign L1[823:820] = sbox[ { round_in[205], state_in[823:820] } ];
	assign L1[819:816] = sbox[ { round_in[204], state_in[819:816] } ];
	assign L1[815:812] = sbox[ { round_in[203], state_in[815:812] } ];
	assign L1[811:808] = sbox[ { round_in[202], state_in[811:808] } ];
	assign L1[807:804] = sbox[ { round_in[201], state_in[807:804] } ];
	assign L1[803:800] = sbox[ { round_in[200], state_in[803:800] } ];
	assign L1[799:796] = sbox[ { round_in[199], state_in[799:796] } ];
	assign L1[795:792] = sbox[ { round_in[198], state_in[795:792] } ];
	assign L1[791:788] = sbox[ { round_in[197], state_in[791:788] } ];
	assign L1[787:784] = sbox[ { round_in[196], state_in[787:784] } ];
	assign L1[783:780] = sbox[ { round_in[195], state_in[783:780] } ];
	assign L1[779:776] = sbox[ { round_in[194], state_in[779:776] } ];
	assign L1[775:772] = sbox[ { round_in[193], state_in[775:772] } ];
	assign L1[771:768] = sbox[ { round_in[192], state_in[771:768] } ];
	assign L1[767:764] = sbox[ { round_in[191], state_in[767:764] } ];
	assign L1[763:760] = sbox[ { round_in[190], state_in[763:760] } ];
	assign L1[759:756] = sbox[ { round_in[189], state_in[759:756] } ];
	assign L1[755:752] = sbox[ { round_in[188], state_in[755:752] } ];
	assign L1[751:748] = sbox[ { round_in[187], state_in[751:748] } ];
	assign L1[747:744] = sbox[ { round_in[186], state_in[747:744] } ];
	assign L1[743:740] = sbox[ { round_in[185], state_in[743:740] } ];
	assign L1[739:736] = sbox[ { round_in[184], state_in[739:736] } ];
	assign L1[735:732] = sbox[ { round_in[183], state_in[735:732] } ];
	assign L1[731:728] = sbox[ { round_in[182], state_in[731:728] } ];
	assign L1[727:724] = sbox[ { round_in[181], state_in[727:724] } ];
	assign L1[723:720] = sbox[ { round_in[180], state_in[723:720] } ];
	assign L1[719:716] = sbox[ { round_in[179], state_in[719:716] } ];
	assign L1[715:712] = sbox[ { round_in[178], state_in[715:712] } ];
	assign L1[711:708] = sbox[ { round_in[177], state_in[711:708] } ];
	assign L1[707:704] = sbox[ { round_in[176], state_in[707:704] } ];
	assign L1[703:700] = sbox[ { round_in[175], state_in[703:700] } ];
	assign L1[699:696] = sbox[ { round_in[174], state_in[699:696] } ];
	assign L1[695:692] = sbox[ { round_in[173], state_in[695:692] } ];
	assign L1[691:688] = sbox[ { round_in[172], state_in[691:688] } ];
	assign L1[687:684] = sbox[ { round_in[171], state_in[687:684] } ];
	assign L1[683:680] = sbox[ { round_in[170], state_in[683:680] } ];
	assign L1[679:676] = sbox[ { round_in[169], state_in[679:676] } ];
	assign L1[675:672] = sbox[ { round_in[168], state_in[675:672] } ];
	assign L1[671:668] = sbox[ { round_in[167], state_in[671:668] } ];
	assign L1[667:664] = sbox[ { round_in[166], state_in[667:664] } ];
	assign L1[663:660] = sbox[ { round_in[165], state_in[663:660] } ];
	assign L1[659:656] = sbox[ { round_in[164], state_in[659:656] } ];
	assign L1[655:652] = sbox[ { round_in[163], state_in[655:652] } ];
	assign L1[651:648] = sbox[ { round_in[162], state_in[651:648] } ];
	assign L1[647:644] = sbox[ { round_in[161], state_in[647:644] } ];
	assign L1[643:640] = sbox[ { round_in[160], state_in[643:640] } ];
	assign L1[639:636] = sbox[ { round_in[159], state_in[639:636] } ];
	assign L1[635:632] = sbox[ { round_in[158], state_in[635:632] } ];
	assign L1[631:628] = sbox[ { round_in[157], state_in[631:628] } ];
	assign L1[627:624] = sbox[ { round_in[156], state_in[627:624] } ];
	assign L1[623:620] = sbox[ { round_in[155], state_in[623:620] } ];
	assign L1[619:616] = sbox[ { round_in[154], state_in[619:616] } ];
	assign L1[615:612] = sbox[ { round_in[153], state_in[615:612] } ];
	assign L1[611:608] = sbox[ { round_in[152], state_in[611:608] } ];
	assign L1[607:604] = sbox[ { round_in[151], state_in[607:604] } ];
	assign L1[603:600] = sbox[ { round_in[150], state_in[603:600] } ];
	assign L1[599:596] = sbox[ { round_in[149], state_in[599:596] } ];
	assign L1[595:592] = sbox[ { round_in[148], state_in[595:592] } ];
	assign L1[591:588] = sbox[ { round_in[147], state_in[591:588] } ];
	assign L1[587:584] = sbox[ { round_in[146], state_in[587:584] } ];
	assign L1[583:580] = sbox[ { round_in[145], state_in[583:580] } ];
	assign L1[579:576] = sbox[ { round_in[144], state_in[579:576] } ];
	assign L1[575:572] = sbox[ { round_in[143], state_in[575:572] } ];
	assign L1[571:568] = sbox[ { round_in[142], state_in[571:568] } ];
	assign L1[567:564] = sbox[ { round_in[141], state_in[567:564] } ];
	assign L1[563:560] = sbox[ { round_in[140], state_in[563:560] } ];
	assign L1[559:556] = sbox[ { round_in[139], state_in[559:556] } ];
	assign L1[555:552] = sbox[ { round_in[138], state_in[555:552] } ];
	assign L1[551:548] = sbox[ { round_in[137], state_in[551:548] } ];
	assign L1[547:544] = sbox[ { round_in[136], state_in[547:544] } ];
	assign L1[543:540] = sbox[ { round_in[135], state_in[543:540] } ];
	assign L1[539:536] = sbox[ { round_in[134], state_in[539:536] } ];
	assign L1[535:532] = sbox[ { round_in[133], state_in[535:532] } ];
	assign L1[531:528] = sbox[ { round_in[132], state_in[531:528] } ];
	assign L1[527:524] = sbox[ { round_in[131], state_in[527:524] } ];
	assign L1[523:520] = sbox[ { round_in[130], state_in[523:520] } ];
	assign L1[519:516] = sbox[ { round_in[129], state_in[519:516] } ];
	assign L1[515:512] = sbox[ { round_in[128], state_in[515:512] } ];
	assign L1[511:508] = sbox[ { round_in[127], state_in[511:508] } ];
	assign L1[507:504] = sbox[ { round_in[126], state_in[507:504] } ];
	assign L1[503:500] = sbox[ { round_in[125], state_in[503:500] } ];
	assign L1[499:496] = sbox[ { round_in[124], state_in[499:496] } ];
	assign L1[495:492] = sbox[ { round_in[123], state_in[495:492] } ];
	assign L1[491:488] = sbox[ { round_in[122], state_in[491:488] } ];
	assign L1[487:484] = sbox[ { round_in[121], state_in[487:484] } ];
	assign L1[483:480] = sbox[ { round_in[120], state_in[483:480] } ];
	assign L1[479:476] = sbox[ { round_in[119], state_in[479:476] } ];
	assign L1[475:472] = sbox[ { round_in[118], state_in[475:472] } ];
	assign L1[471:468] = sbox[ { round_in[117], state_in[471:468] } ];
	assign L1[467:464] = sbox[ { round_in[116], state_in[467:464] } ];
	assign L1[463:460] = sbox[ { round_in[115], state_in[463:460] } ];
	assign L1[459:456] = sbox[ { round_in[114], state_in[459:456] } ];
	assign L1[455:452] = sbox[ { round_in[113], state_in[455:452] } ];
	assign L1[451:448] = sbox[ { round_in[112], state_in[451:448] } ];
	assign L1[447:444] = sbox[ { round_in[111], state_in[447:444] } ];
	assign L1[443:440] = sbox[ { round_in[110], state_in[443:440] } ];
	assign L1[439:436] = sbox[ { round_in[109], state_in[439:436] } ];
	assign L1[435:432] = sbox[ { round_in[108], state_in[435:432] } ];
	assign L1[431:428] = sbox[ { round_in[107], state_in[431:428] } ];
	assign L1[427:424] = sbox[ { round_in[106], state_in[427:424] } ];
	assign L1[423:420] = sbox[ { round_in[105], state_in[423:420] } ];
	assign L1[419:416] = sbox[ { round_in[104], state_in[419:416] } ];
	assign L1[415:412] = sbox[ { round_in[103], state_in[415:412] } ];
	assign L1[411:408] = sbox[ { round_in[102], state_in[411:408] } ];
	assign L1[407:404] = sbox[ { round_in[101], state_in[407:404] } ];
	assign L1[403:400] = sbox[ { round_in[100], state_in[403:400] } ];
	assign L1[399:396] = sbox[ { round_in[99], state_in[399:396] } ];
	assign L1[395:392] = sbox[ { round_in[98], state_in[395:392] } ];
	assign L1[391:388] = sbox[ { round_in[97], state_in[391:388] } ];
	assign L1[387:384] = sbox[ { round_in[96], state_in[387:384] } ];
	assign L1[383:380] = sbox[ { round_in[95], state_in[383:380] } ];
	assign L1[379:376] = sbox[ { round_in[94], state_in[379:376] } ];
	assign L1[375:372] = sbox[ { round_in[93], state_in[375:372] } ];
	assign L1[371:368] = sbox[ { round_in[92], state_in[371:368] } ];
	assign L1[367:364] = sbox[ { round_in[91], state_in[367:364] } ];
	assign L1[363:360] = sbox[ { round_in[90], state_in[363:360] } ];
	assign L1[359:356] = sbox[ { round_in[89], state_in[359:356] } ];
	assign L1[355:352] = sbox[ { round_in[88], state_in[355:352] } ];
	assign L1[351:348] = sbox[ { round_in[87], state_in[351:348] } ];
	assign L1[347:344] = sbox[ { round_in[86], state_in[347:344] } ];
	assign L1[343:340] = sbox[ { round_in[85], state_in[343:340] } ];
	assign L1[339:336] = sbox[ { round_in[84], state_in[339:336] } ];
	assign L1[335:332] = sbox[ { round_in[83], state_in[335:332] } ];
	assign L1[331:328] = sbox[ { round_in[82], state_in[331:328] } ];
	assign L1[327:324] = sbox[ { round_in[81], state_in[327:324] } ];
	assign L1[323:320] = sbox[ { round_in[80], state_in[323:320] } ];
	assign L1[319:316] = sbox[ { round_in[79], state_in[319:316] } ];
	assign L1[315:312] = sbox[ { round_in[78], state_in[315:312] } ];
	assign L1[311:308] = sbox[ { round_in[77], state_in[311:308] } ];
	assign L1[307:304] = sbox[ { round_in[76], state_in[307:304] } ];
	assign L1[303:300] = sbox[ { round_in[75], state_in[303:300] } ];
	assign L1[299:296] = sbox[ { round_in[74], state_in[299:296] } ];
	assign L1[295:292] = sbox[ { round_in[73], state_in[295:292] } ];
	assign L1[291:288] = sbox[ { round_in[72], state_in[291:288] } ];
	assign L1[287:284] = sbox[ { round_in[71], state_in[287:284] } ];
	assign L1[283:280] = sbox[ { round_in[70], state_in[283:280] } ];
	assign L1[279:276] = sbox[ { round_in[69], state_in[279:276] } ];
	assign L1[275:272] = sbox[ { round_in[68], state_in[275:272] } ];
	assign L1[271:268] = sbox[ { round_in[67], state_in[271:268] } ];
	assign L1[267:264] = sbox[ { round_in[66], state_in[267:264] } ];
	assign L1[263:260] = sbox[ { round_in[65], state_in[263:260] } ];
	assign L1[259:256] = sbox[ { round_in[64], state_in[259:256] } ];
	assign L1[255:252] = sbox[ { round_in[63], state_in[255:252] } ];
	assign L1[251:248] = sbox[ { round_in[62], state_in[251:248] } ];
	assign L1[247:244] = sbox[ { round_in[61], state_in[247:244] } ];
	assign L1[243:240] = sbox[ { round_in[60], state_in[243:240] } ];
	assign L1[239:236] = sbox[ { round_in[59], state_in[239:236] } ];
	assign L1[235:232] = sbox[ { round_in[58], state_in[235:232] } ];
	assign L1[231:228] = sbox[ { round_in[57], state_in[231:228] } ];
	assign L1[227:224] = sbox[ { round_in[56], state_in[227:224] } ];
	assign L1[223:220] = sbox[ { round_in[55], state_in[223:220] } ];
	assign L1[219:216] = sbox[ { round_in[54], state_in[219:216] } ];
	assign L1[215:212] = sbox[ { round_in[53], state_in[215:212] } ];
	assign L1[211:208] = sbox[ { round_in[52], state_in[211:208] } ];
	assign L1[207:204] = sbox[ { round_in[51], state_in[207:204] } ];
	assign L1[203:200] = sbox[ { round_in[50], state_in[203:200] } ];
	assign L1[199:196] = sbox[ { round_in[49], state_in[199:196] } ];
	assign L1[195:192] = sbox[ { round_in[48], state_in[195:192] } ];
	assign L1[191:188] = sbox[ { round_in[47], state_in[191:188] } ];
	assign L1[187:184] = sbox[ { round_in[46], state_in[187:184] } ];
	assign L1[183:180] = sbox[ { round_in[45], state_in[183:180] } ];
	assign L1[179:176] = sbox[ { round_in[44], state_in[179:176] } ];
	assign L1[175:172] = sbox[ { round_in[43], state_in[175:172] } ];
	assign L1[171:168] = sbox[ { round_in[42], state_in[171:168] } ];
	assign L1[167:164] = sbox[ { round_in[41], state_in[167:164] } ];
	assign L1[163:160] = sbox[ { round_in[40], state_in[163:160] } ];
	assign L1[159:156] = sbox[ { round_in[39], state_in[159:156] } ];
	assign L1[155:152] = sbox[ { round_in[38], state_in[155:152] } ];
	assign L1[151:148] = sbox[ { round_in[37], state_in[151:148] } ];
	assign L1[147:144] = sbox[ { round_in[36], state_in[147:144] } ];
	assign L1[143:140] = sbox[ { round_in[35], state_in[143:140] } ];
	assign L1[139:136] = sbox[ { round_in[34], state_in[139:136] } ];
	assign L1[135:132] = sbox[ { round_in[33], state_in[135:132] } ];
	assign L1[131:128] = sbox[ { round_in[32], state_in[131:128] } ];
	assign L1[127:124] = sbox[ { round_in[31], state_in[127:124] } ];
	assign L1[123:120] = sbox[ { round_in[30], state_in[123:120] } ];
	assign L1[119:116] = sbox[ { round_in[29], state_in[119:116] } ];
	assign L1[115:112] = sbox[ { round_in[28], state_in[115:112] } ];
	assign L1[111:108] = sbox[ { round_in[27], state_in[111:108] } ];
	assign L1[107:104] = sbox[ { round_in[26], state_in[107:104] } ];
	assign L1[103:100] = sbox[ { round_in[25], state_in[103:100] } ];
	assign L1[99:96] = sbox[ { round_in[24], state_in[99:96] } ];
	assign L1[95:92] = sbox[ { round_in[23], state_in[95:92] } ];
	assign L1[91:88] = sbox[ { round_in[22], state_in[91:88] } ];
	assign L1[87:84] = sbox[ { round_in[21], state_in[87:84] } ];
	assign L1[83:80] = sbox[ { round_in[20], state_in[83:80] } ];
	assign L1[79:76] = sbox[ { round_in[19], state_in[79:76] } ];
	assign L1[75:72] = sbox[ { round_in[18], state_in[75:72] } ];
	assign L1[71:68] = sbox[ { round_in[17], state_in[71:68] } ];
	assign L1[67:64] = sbox[ { round_in[16], state_in[67:64] } ];
	assign L1[63:60] = sbox[ { round_in[15], state_in[63:60] } ];
	assign L1[59:56] = sbox[ { round_in[14], state_in[59:56] } ];
	assign L1[55:52] = sbox[ { round_in[13], state_in[55:52] } ];
	assign L1[51:48] = sbox[ { round_in[12], state_in[51:48] } ];
	assign L1[47:44] = sbox[ { round_in[11], state_in[47:44] } ];
	assign L1[43:40] = sbox[ { round_in[10], state_in[43:40] } ];
	assign L1[39:36] = sbox[ { round_in[9], state_in[39:36] } ];
	assign L1[35:32] = sbox[ { round_in[8], state_in[35:32] } ];
	assign L1[31:28] = sbox[ { round_in[7], state_in[31:28] } ];
	assign L1[27:24] = sbox[ { round_in[6], state_in[27:24] } ];
	assign L1[23:20] = sbox[ { round_in[5], state_in[23:20] } ];
	assign L1[19:16] = sbox[ { round_in[4], state_in[19:16] } ];
	assign L1[15:12] = sbox[ { round_in[3], state_in[15:12] } ];
	assign L1[11:8] = sbox[ { round_in[2], state_in[11:8] } ];
	assign L1[7:4] = sbox[ { round_in[1], state_in[7:4] } ];
	assign L1[3:0] = sbox[ { round_in[0], state_in[3:0] } ];

	assign out[1023:1020] = { L1[1015]^L1[1010], L1[1014]^L1[1009], L1[1013]^L1[1008]^L1[1011], L1[1012]^L1[1011] };
	assign out[1019:1016] = { L1[1019]^L1[1022]^L1[1017], L1[1018]^L1[1021]^L1[1016]^L1[1019], L1[1017]^L1[1020]^L1[1019]^L1[1023]^L1[1018], L1[1016]^L1[1023]^L1[1018] };
	assign out[1015:1012] = { L1[999]^L1[994], L1[998]^L1[993], L1[997]^L1[992]^L1[995], L1[996]^L1[995] };
	assign out[1011:1008] = { L1[1003]^L1[1006]^L1[1001], L1[1002]^L1[1005]^L1[1000]^L1[1003], L1[1001]^L1[1004]^L1[1003]^L1[1007]^L1[1002], L1[1000]^L1[1007]^L1[1002] };
	assign out[1007:1004] = { L1[983]^L1[978], L1[982]^L1[977], L1[981]^L1[976]^L1[979], L1[980]^L1[979] };
	assign out[1003:1000] = { L1[987]^L1[990]^L1[985], L1[986]^L1[989]^L1[984]^L1[987], L1[985]^L1[988]^L1[987]^L1[991]^L1[986], L1[984]^L1[991]^L1[986] };
	assign out[999:996]   = { L1[967]^L1[962], L1[966]^L1[961], L1[965]^L1[960]^L1[963], L1[964]^L1[963] };
	assign out[995:992]   = { L1[971]^L1[974]^L1[969], L1[970]^L1[973]^L1[968]^L1[971], L1[969]^L1[972]^L1[971]^L1[975]^L1[970], L1[968]^L1[975]^L1[970] };
	assign out[991:988]   = { L1[951]^L1[946], L1[950]^L1[945], L1[949]^L1[944]^L1[947], L1[948]^L1[947] };
	assign out[987:984]   = { L1[955]^L1[958]^L1[953], L1[954]^L1[957]^L1[952]^L1[955], L1[953]^L1[956]^L1[955]^L1[959]^L1[954], L1[952]^L1[959]^L1[954] };
	assign out[983:980]   = { L1[935]^L1[930], L1[934]^L1[929], L1[933]^L1[928]^L1[931], L1[932]^L1[931] };
	assign out[979:976]   = { L1[939]^L1[942]^L1[937], L1[938]^L1[941]^L1[936]^L1[939], L1[937]^L1[940]^L1[939]^L1[943]^L1[938], L1[936]^L1[943]^L1[938] };
	assign out[975:972]   = { L1[919]^L1[914], L1[918]^L1[913], L1[917]^L1[912]^L1[915], L1[916]^L1[915] };
	assign out[971:968]   = { L1[923]^L1[926]^L1[921], L1[922]^L1[925]^L1[920]^L1[923], L1[921]^L1[924]^L1[923]^L1[927]^L1[922], L1[920]^L1[927]^L1[922] };
	assign out[967:964]   = { L1[903]^L1[898], L1[902]^L1[897], L1[901]^L1[896]^L1[899], L1[900]^L1[899] };
	assign out[963:960]   = { L1[907]^L1[910]^L1[905], L1[906]^L1[909]^L1[904]^L1[907], L1[905]^L1[908]^L1[907]^L1[911]^L1[906], L1[904]^L1[911]^L1[906] };
	assign out[959:956]   = { L1[887]^L1[882], L1[886]^L1[881], L1[885]^L1[880]^L1[883], L1[884]^L1[883] };
	assign out[955:952]   = { L1[891]^L1[894]^L1[889], L1[890]^L1[893]^L1[888]^L1[891], L1[889]^L1[892]^L1[891]^L1[895]^L1[890], L1[888]^L1[895]^L1[890] };
	assign out[951:948]   = { L1[871]^L1[866], L1[870]^L1[865], L1[869]^L1[864]^L1[867], L1[868]^L1[867] };
	assign out[947:944]   = { L1[875]^L1[878]^L1[873], L1[874]^L1[877]^L1[872]^L1[875], L1[873]^L1[876]^L1[875]^L1[879]^L1[874], L1[872]^L1[879]^L1[874] };
	assign out[943:940]   = { L1[855]^L1[850], L1[854]^L1[849], L1[853]^L1[848]^L1[851], L1[852]^L1[851] };
	assign out[939:936]   = { L1[859]^L1[862]^L1[857], L1[858]^L1[861]^L1[856]^L1[859], L1[857]^L1[860]^L1[859]^L1[863]^L1[858], L1[856]^L1[863]^L1[858] };
	assign out[935:932]   = { L1[839]^L1[834], L1[838]^L1[833], L1[837]^L1[832]^L1[835], L1[836]^L1[835] };
	assign out[931:928]   = { L1[843]^L1[846]^L1[841], L1[842]^L1[845]^L1[840]^L1[843], L1[841]^L1[844]^L1[843]^L1[847]^L1[842], L1[840]^L1[847]^L1[842] };
	assign out[927:924]   = { L1[823]^L1[818], L1[822]^L1[817], L1[821]^L1[816]^L1[819], L1[820]^L1[819] };
	assign out[923:920]   = { L1[827]^L1[830]^L1[825], L1[826]^L1[829]^L1[824]^L1[827], L1[825]^L1[828]^L1[827]^L1[831]^L1[826], L1[824]^L1[831]^L1[826] };
	assign out[919:916]   = { L1[807]^L1[802], L1[806]^L1[801], L1[805]^L1[800]^L1[803], L1[804]^L1[803] };
	assign out[915:912]   = { L1[811]^L1[814]^L1[809], L1[810]^L1[813]^L1[808]^L1[811], L1[809]^L1[812]^L1[811]^L1[815]^L1[810], L1[808]^L1[815]^L1[810] };
	assign out[911:908]   = { L1[791]^L1[786], L1[790]^L1[785], L1[789]^L1[784]^L1[787], L1[788]^L1[787] };
	assign out[907:904]   = { L1[795]^L1[798]^L1[793], L1[794]^L1[797]^L1[792]^L1[795], L1[793]^L1[796]^L1[795]^L1[799]^L1[794], L1[792]^L1[799]^L1[794] };
	assign out[903:900]   = { L1[775]^L1[770], L1[774]^L1[769], L1[773]^L1[768]^L1[771], L1[772]^L1[771] };
	assign out[899:896]   = { L1[779]^L1[782]^L1[777], L1[778]^L1[781]^L1[776]^L1[779], L1[777]^L1[780]^L1[779]^L1[783]^L1[778], L1[776]^L1[783]^L1[778] };
	assign out[895:892]   = { L1[759]^L1[754], L1[758]^L1[753], L1[757]^L1[752]^L1[755], L1[756]^L1[755] };
	assign out[891:888]   = { L1[763]^L1[766]^L1[761], L1[762]^L1[765]^L1[760]^L1[763], L1[761]^L1[764]^L1[763]^L1[767]^L1[762], L1[760]^L1[767]^L1[762] };
	assign out[887:884]   = { L1[743]^L1[738], L1[742]^L1[737], L1[741]^L1[736]^L1[739], L1[740]^L1[739] };
	assign out[883:880]   = { L1[747]^L1[750]^L1[745], L1[746]^L1[749]^L1[744]^L1[747], L1[745]^L1[748]^L1[747]^L1[751]^L1[746], L1[744]^L1[751]^L1[746] };
	assign out[879:876]   = { L1[727]^L1[722], L1[726]^L1[721], L1[725]^L1[720]^L1[723], L1[724]^L1[723] };
	assign out[875:872]   = { L1[731]^L1[734]^L1[729], L1[730]^L1[733]^L1[728]^L1[731], L1[729]^L1[732]^L1[731]^L1[735]^L1[730], L1[728]^L1[735]^L1[730] };
	assign out[871:868]   = { L1[711]^L1[706], L1[710]^L1[705], L1[709]^L1[704]^L1[707], L1[708]^L1[707] };
	assign out[867:864]   = { L1[715]^L1[718]^L1[713], L1[714]^L1[717]^L1[712]^L1[715], L1[713]^L1[716]^L1[715]^L1[719]^L1[714], L1[712]^L1[719]^L1[714] };
	assign out[863:860]   = { L1[695]^L1[690], L1[694]^L1[689], L1[693]^L1[688]^L1[691], L1[692]^L1[691] };
	assign out[859:856]   = { L1[699]^L1[702]^L1[697], L1[698]^L1[701]^L1[696]^L1[699], L1[697]^L1[700]^L1[699]^L1[703]^L1[698], L1[696]^L1[703]^L1[698] };
	assign out[855:852]   = { L1[679]^L1[674], L1[678]^L1[673], L1[677]^L1[672]^L1[675], L1[676]^L1[675] };
	assign out[851:848]   = { L1[683]^L1[686]^L1[681], L1[682]^L1[685]^L1[680]^L1[683], L1[681]^L1[684]^L1[683]^L1[687]^L1[682], L1[680]^L1[687]^L1[682] };
	assign out[847:844]   = { L1[663]^L1[658], L1[662]^L1[657], L1[661]^L1[656]^L1[659], L1[660]^L1[659] };
	assign out[843:840]   = { L1[667]^L1[670]^L1[665], L1[666]^L1[669]^L1[664]^L1[667], L1[665]^L1[668]^L1[667]^L1[671]^L1[666], L1[664]^L1[671]^L1[666] };
	assign out[839:836]   = { L1[647]^L1[642], L1[646]^L1[641], L1[645]^L1[640]^L1[643], L1[644]^L1[643] };
	assign out[835:832]   = { L1[651]^L1[654]^L1[649], L1[650]^L1[653]^L1[648]^L1[651], L1[649]^L1[652]^L1[651]^L1[655]^L1[650], L1[648]^L1[655]^L1[650] };
	assign out[831:828]   = { L1[631]^L1[626], L1[630]^L1[625], L1[629]^L1[624]^L1[627], L1[628]^L1[627] };
	assign out[827:824]   = { L1[635]^L1[638]^L1[633], L1[634]^L1[637]^L1[632]^L1[635], L1[633]^L1[636]^L1[635]^L1[639]^L1[634], L1[632]^L1[639]^L1[634] };
	assign out[823:820]   = { L1[615]^L1[610], L1[614]^L1[609], L1[613]^L1[608]^L1[611], L1[612]^L1[611] };
	assign out[819:816]   = { L1[619]^L1[622]^L1[617], L1[618]^L1[621]^L1[616]^L1[619], L1[617]^L1[620]^L1[619]^L1[623]^L1[618], L1[616]^L1[623]^L1[618] };
	assign out[815:812]   = { L1[599]^L1[594], L1[598]^L1[593], L1[597]^L1[592]^L1[595], L1[596]^L1[595] };
	assign out[811:808]   = { L1[603]^L1[606]^L1[601], L1[602]^L1[605]^L1[600]^L1[603], L1[601]^L1[604]^L1[603]^L1[607]^L1[602], L1[600]^L1[607]^L1[602] };
	assign out[807:804]   = { L1[583]^L1[578], L1[582]^L1[577], L1[581]^L1[576]^L1[579], L1[580]^L1[579] };
	assign out[803:800]   = { L1[587]^L1[590]^L1[585], L1[586]^L1[589]^L1[584]^L1[587], L1[585]^L1[588]^L1[587]^L1[591]^L1[586], L1[584]^L1[591]^L1[586] };
	assign out[799:796]   = { L1[567]^L1[562], L1[566]^L1[561], L1[565]^L1[560]^L1[563], L1[564]^L1[563] };
	assign out[795:792]   = { L1[571]^L1[574]^L1[569], L1[570]^L1[573]^L1[568]^L1[571], L1[569]^L1[572]^L1[571]^L1[575]^L1[570], L1[568]^L1[575]^L1[570] };
	assign out[791:788]   = { L1[551]^L1[546], L1[550]^L1[545], L1[549]^L1[544]^L1[547], L1[548]^L1[547] };
	assign out[787:784]   = { L1[555]^L1[558]^L1[553], L1[554]^L1[557]^L1[552]^L1[555], L1[553]^L1[556]^L1[555]^L1[559]^L1[554], L1[552]^L1[559]^L1[554] };
	assign out[783:780]   = { L1[535]^L1[530], L1[534]^L1[529], L1[533]^L1[528]^L1[531], L1[532]^L1[531] };
	assign out[779:776]   = { L1[539]^L1[542]^L1[537], L1[538]^L1[541]^L1[536]^L1[539], L1[537]^L1[540]^L1[539]^L1[543]^L1[538], L1[536]^L1[543]^L1[538] };
	assign out[775:772]   = { L1[519]^L1[514], L1[518]^L1[513], L1[517]^L1[512]^L1[515], L1[516]^L1[515] };
	assign out[771:768]   = { L1[523]^L1[526]^L1[521], L1[522]^L1[525]^L1[520]^L1[523], L1[521]^L1[524]^L1[523]^L1[527]^L1[522], L1[520]^L1[527]^L1[522] };
	assign out[767:764]   = { L1[503]^L1[498], L1[502]^L1[497], L1[501]^L1[496]^L1[499], L1[500]^L1[499] };
	assign out[763:760]   = { L1[507]^L1[510]^L1[505], L1[506]^L1[509]^L1[504]^L1[507], L1[505]^L1[508]^L1[507]^L1[511]^L1[506], L1[504]^L1[511]^L1[506] };
	assign out[759:756]   = { L1[487]^L1[482], L1[486]^L1[481], L1[485]^L1[480]^L1[483], L1[484]^L1[483] };
	assign out[755:752]   = { L1[491]^L1[494]^L1[489], L1[490]^L1[493]^L1[488]^L1[491], L1[489]^L1[492]^L1[491]^L1[495]^L1[490], L1[488]^L1[495]^L1[490] };
	assign out[751:748]   = { L1[471]^L1[466], L1[470]^L1[465], L1[469]^L1[464]^L1[467], L1[468]^L1[467] };
	assign out[747:744]   = { L1[475]^L1[478]^L1[473], L1[474]^L1[477]^L1[472]^L1[475], L1[473]^L1[476]^L1[475]^L1[479]^L1[474], L1[472]^L1[479]^L1[474] };
	assign out[743:740]   = { L1[455]^L1[450], L1[454]^L1[449], L1[453]^L1[448]^L1[451], L1[452]^L1[451] };
	assign out[739:736]   = { L1[459]^L1[462]^L1[457], L1[458]^L1[461]^L1[456]^L1[459], L1[457]^L1[460]^L1[459]^L1[463]^L1[458], L1[456]^L1[463]^L1[458] };
	assign out[735:732]   = { L1[439]^L1[434], L1[438]^L1[433], L1[437]^L1[432]^L1[435], L1[436]^L1[435] };
	assign out[731:728]   = { L1[443]^L1[446]^L1[441], L1[442]^L1[445]^L1[440]^L1[443], L1[441]^L1[444]^L1[443]^L1[447]^L1[442], L1[440]^L1[447]^L1[442] };
	assign out[727:724]   = { L1[423]^L1[418], L1[422]^L1[417], L1[421]^L1[416]^L1[419], L1[420]^L1[419] };
	assign out[723:720]   = { L1[427]^L1[430]^L1[425], L1[426]^L1[429]^L1[424]^L1[427], L1[425]^L1[428]^L1[427]^L1[431]^L1[426], L1[424]^L1[431]^L1[426] };
	assign out[719:716]   = { L1[407]^L1[402], L1[406]^L1[401], L1[405]^L1[400]^L1[403], L1[404]^L1[403] };
	assign out[715:712]   = { L1[411]^L1[414]^L1[409], L1[410]^L1[413]^L1[408]^L1[411], L1[409]^L1[412]^L1[411]^L1[415]^L1[410], L1[408]^L1[415]^L1[410] };
	assign out[711:708]   = { L1[391]^L1[386], L1[390]^L1[385], L1[389]^L1[384]^L1[387], L1[388]^L1[387] };
	assign out[707:704]   = { L1[395]^L1[398]^L1[393], L1[394]^L1[397]^L1[392]^L1[395], L1[393]^L1[396]^L1[395]^L1[399]^L1[394], L1[392]^L1[399]^L1[394] };
	assign out[703:700]   = { L1[375]^L1[370], L1[374]^L1[369], L1[373]^L1[368]^L1[371], L1[372]^L1[371] };
	assign out[699:696]   = { L1[379]^L1[382]^L1[377], L1[378]^L1[381]^L1[376]^L1[379], L1[377]^L1[380]^L1[379]^L1[383]^L1[378], L1[376]^L1[383]^L1[378] };
	assign out[695:692]   = { L1[359]^L1[354], L1[358]^L1[353], L1[357]^L1[352]^L1[355], L1[356]^L1[355] };
	assign out[691:688]   = { L1[363]^L1[366]^L1[361], L1[362]^L1[365]^L1[360]^L1[363], L1[361]^L1[364]^L1[363]^L1[367]^L1[362], L1[360]^L1[367]^L1[362] };
	assign out[687:684]   = { L1[343]^L1[338], L1[342]^L1[337], L1[341]^L1[336]^L1[339], L1[340]^L1[339] };
	assign out[683:680]   = { L1[347]^L1[350]^L1[345], L1[346]^L1[349]^L1[344]^L1[347], L1[345]^L1[348]^L1[347]^L1[351]^L1[346], L1[344]^L1[351]^L1[346] };
	assign out[679:676]   = { L1[327]^L1[322], L1[326]^L1[321], L1[325]^L1[320]^L1[323], L1[324]^L1[323] };
	assign out[675:672]   = { L1[331]^L1[334]^L1[329], L1[330]^L1[333]^L1[328]^L1[331], L1[329]^L1[332]^L1[331]^L1[335]^L1[330], L1[328]^L1[335]^L1[330] };
	assign out[671:668]   = { L1[311]^L1[306], L1[310]^L1[305], L1[309]^L1[304]^L1[307], L1[308]^L1[307] };
	assign out[667:664]   = { L1[315]^L1[318]^L1[313], L1[314]^L1[317]^L1[312]^L1[315], L1[313]^L1[316]^L1[315]^L1[319]^L1[314], L1[312]^L1[319]^L1[314] };
	assign out[663:660]   = { L1[295]^L1[290], L1[294]^L1[289], L1[293]^L1[288]^L1[291], L1[292]^L1[291] };
	assign out[659:656]   = { L1[299]^L1[302]^L1[297], L1[298]^L1[301]^L1[296]^L1[299], L1[297]^L1[300]^L1[299]^L1[303]^L1[298], L1[296]^L1[303]^L1[298] };
	assign out[655:652]   = { L1[279]^L1[274], L1[278]^L1[273], L1[277]^L1[272]^L1[275], L1[276]^L1[275] };
	assign out[651:648]   = { L1[283]^L1[286]^L1[281], L1[282]^L1[285]^L1[280]^L1[283], L1[281]^L1[284]^L1[283]^L1[287]^L1[282], L1[280]^L1[287]^L1[282] };
	assign out[647:644]   = { L1[263]^L1[258], L1[262]^L1[257], L1[261]^L1[256]^L1[259], L1[260]^L1[259] };
	assign out[643:640]   = { L1[267]^L1[270]^L1[265], L1[266]^L1[269]^L1[264]^L1[267], L1[265]^L1[268]^L1[267]^L1[271]^L1[266], L1[264]^L1[271]^L1[266] };
	assign out[639:636]   = { L1[247]^L1[242], L1[246]^L1[241], L1[245]^L1[240]^L1[243], L1[244]^L1[243] };
	assign out[635:632]   = { L1[251]^L1[254]^L1[249], L1[250]^L1[253]^L1[248]^L1[251], L1[249]^L1[252]^L1[251]^L1[255]^L1[250], L1[248]^L1[255]^L1[250] };
	assign out[631:628]   = { L1[231]^L1[226], L1[230]^L1[225], L1[229]^L1[224]^L1[227], L1[228]^L1[227] };
	assign out[627:624]   = { L1[235]^L1[238]^L1[233], L1[234]^L1[237]^L1[232]^L1[235], L1[233]^L1[236]^L1[235]^L1[239]^L1[234], L1[232]^L1[239]^L1[234] };
	assign out[623:620]   = { L1[215]^L1[210], L1[214]^L1[209], L1[213]^L1[208]^L1[211], L1[212]^L1[211] };
	assign out[619:616]   = { L1[219]^L1[222]^L1[217], L1[218]^L1[221]^L1[216]^L1[219], L1[217]^L1[220]^L1[219]^L1[223]^L1[218], L1[216]^L1[223]^L1[218] };
	assign out[615:612]   = { L1[199]^L1[194], L1[198]^L1[193], L1[197]^L1[192]^L1[195], L1[196]^L1[195] };
	assign out[611:608]   = { L1[203]^L1[206]^L1[201], L1[202]^L1[205]^L1[200]^L1[203], L1[201]^L1[204]^L1[203]^L1[207]^L1[202], L1[200]^L1[207]^L1[202] };
	assign out[607:604]   = { L1[183]^L1[178], L1[182]^L1[177], L1[181]^L1[176]^L1[179], L1[180]^L1[179] };
	assign out[603:600]   = { L1[187]^L1[190]^L1[185], L1[186]^L1[189]^L1[184]^L1[187], L1[185]^L1[188]^L1[187]^L1[191]^L1[186], L1[184]^L1[191]^L1[186] };
	assign out[599:596]   = { L1[167]^L1[162], L1[166]^L1[161], L1[165]^L1[160]^L1[163], L1[164]^L1[163] };
	assign out[595:592]   = { L1[171]^L1[174]^L1[169], L1[170]^L1[173]^L1[168]^L1[171], L1[169]^L1[172]^L1[171]^L1[175]^L1[170], L1[168]^L1[175]^L1[170] };
	assign out[591:588]   = { L1[151]^L1[146], L1[150]^L1[145], L1[149]^L1[144]^L1[147], L1[148]^L1[147] };
	assign out[587:584]   = { L1[155]^L1[158]^L1[153], L1[154]^L1[157]^L1[152]^L1[155], L1[153]^L1[156]^L1[155]^L1[159]^L1[154], L1[152]^L1[159]^L1[154] };
	assign out[583:580]   = { L1[135]^L1[130], L1[134]^L1[129], L1[133]^L1[128]^L1[131], L1[132]^L1[131] };
	assign out[579:576]   = { L1[139]^L1[142]^L1[137], L1[138]^L1[141]^L1[136]^L1[139], L1[137]^L1[140]^L1[139]^L1[143]^L1[138], L1[136]^L1[143]^L1[138] };
	assign out[575:572]   = { L1[119]^L1[114], L1[118]^L1[113], L1[117]^L1[112]^L1[115], L1[116]^L1[115] };
	assign out[571:568]   = { L1[123]^L1[126]^L1[121], L1[122]^L1[125]^L1[120]^L1[123], L1[121]^L1[124]^L1[123]^L1[127]^L1[122], L1[120]^L1[127]^L1[122] };
	assign out[567:564]   = { L1[103]^L1[98], L1[102]^L1[97], L1[101]^L1[96]^L1[99], L1[100]^L1[99] };
	assign out[563:560]   = { L1[107]^L1[110]^L1[105], L1[106]^L1[109]^L1[104]^L1[107], L1[105]^L1[108]^L1[107]^L1[111]^L1[106], L1[104]^L1[111]^L1[106] };
	assign out[559:556]   = { L1[87]^L1[82], L1[86]^L1[81], L1[85]^L1[80]^L1[83], L1[84]^L1[83] };
	assign out[555:552]   = { L1[91]^L1[94]^L1[89], L1[90]^L1[93]^L1[88]^L1[91], L1[89]^L1[92]^L1[91]^L1[95]^L1[90], L1[88]^L1[95]^L1[90] };
	assign out[551:548]   = { L1[71]^L1[66], L1[70]^L1[65], L1[69]^L1[64]^L1[67], L1[68]^L1[67] };
	assign out[547:544]   = { L1[75]^L1[78]^L1[73], L1[74]^L1[77]^L1[72]^L1[75], L1[73]^L1[76]^L1[75]^L1[79]^L1[74], L1[72]^L1[79]^L1[74] };
	assign out[543:540]   = { L1[55]^L1[50], L1[54]^L1[49], L1[53]^L1[48]^L1[51], L1[52]^L1[51] };
	assign out[539:536]   = { L1[59]^L1[62]^L1[57], L1[58]^L1[61]^L1[56]^L1[59], L1[57]^L1[60]^L1[59]^L1[63]^L1[58], L1[56]^L1[63]^L1[58] };
	assign out[535:532]   = { L1[39]^L1[34], L1[38]^L1[33], L1[37]^L1[32]^L1[35], L1[36]^L1[35] };
	assign out[531:528]   = { L1[43]^L1[46]^L1[41], L1[42]^L1[45]^L1[40]^L1[43], L1[41]^L1[44]^L1[43]^L1[47]^L1[42], L1[40]^L1[47]^L1[42] };
	assign out[527:524]   = { L1[23]^L1[18], L1[22]^L1[17], L1[21]^L1[16]^L1[19], L1[20]^L1[19] };
	assign out[523:520]   = { L1[27]^L1[30]^L1[25], L1[26]^L1[29]^L1[24]^L1[27], L1[25]^L1[28]^L1[27]^L1[31]^L1[26], L1[24]^L1[31]^L1[26] };
	assign out[519:516]   = { L1[7]^L1[2], L1[6]^L1[1], L1[5]^L1[0]^L1[3], L1[4]^L1[3] };
	assign out[515:512]   = { L1[11]^L1[14]^L1[9], L1[10]^L1[13]^L1[8]^L1[11], L1[9]^L1[12]^L1[11]^L1[15]^L1[10], L1[8]^L1[15]^L1[10] };
	assign out[511:508]   = { L1[1023]^L1[1018], L1[1022]^L1[1017], L1[1021]^L1[1016]^L1[1019], L1[1020]^L1[1019] };
	assign out[507:504]   = { L1[1011]^L1[1014]^L1[1009], L1[1010]^L1[1013]^L1[1008]^L1[1011], L1[1009]^L1[1012]^L1[1011]^L1[1015]^L1[1010], L1[1008]^L1[1015]^L1[1010] };
	assign out[503:500]   = { L1[1007]^L1[1002], L1[1006]^L1[1001], L1[1005]^L1[1000]^L1[1003], L1[1004]^L1[1003] };
	assign out[499:496]   = { L1[995]^L1[998]^L1[993], L1[994]^L1[997]^L1[992]^L1[995], L1[993]^L1[996]^L1[995]^L1[999]^L1[994], L1[992]^L1[999]^L1[994] };
	assign out[495:492]   = { L1[991]^L1[986], L1[990]^L1[985], L1[989]^L1[984]^L1[987], L1[988]^L1[987] };
	assign out[491:488]   = { L1[979]^L1[982]^L1[977], L1[978]^L1[981]^L1[976]^L1[979], L1[977]^L1[980]^L1[979]^L1[983]^L1[978], L1[976]^L1[983]^L1[978] };
	assign out[487:484]   = { L1[975]^L1[970], L1[974]^L1[969], L1[973]^L1[968]^L1[971], L1[972]^L1[971] };
	assign out[483:480]   = { L1[963]^L1[966]^L1[961], L1[962]^L1[965]^L1[960]^L1[963], L1[961]^L1[964]^L1[963]^L1[967]^L1[962], L1[960]^L1[967]^L1[962] };
	assign out[479:476]   = { L1[959]^L1[954], L1[958]^L1[953], L1[957]^L1[952]^L1[955], L1[956]^L1[955] };
	assign out[475:472]   = { L1[947]^L1[950]^L1[945], L1[946]^L1[949]^L1[944]^L1[947], L1[945]^L1[948]^L1[947]^L1[951]^L1[946], L1[944]^L1[951]^L1[946] };
	assign out[471:468]   = { L1[943]^L1[938], L1[942]^L1[937], L1[941]^L1[936]^L1[939], L1[940]^L1[939] };
	assign out[467:464]   = { L1[931]^L1[934]^L1[929], L1[930]^L1[933]^L1[928]^L1[931], L1[929]^L1[932]^L1[931]^L1[935]^L1[930], L1[928]^L1[935]^L1[930] };
	assign out[463:460]   = { L1[927]^L1[922], L1[926]^L1[921], L1[925]^L1[920]^L1[923], L1[924]^L1[923] };
	assign out[459:456]   = { L1[915]^L1[918]^L1[913], L1[914]^L1[917]^L1[912]^L1[915], L1[913]^L1[916]^L1[915]^L1[919]^L1[914], L1[912]^L1[919]^L1[914] };
	assign out[455:452]   = { L1[911]^L1[906], L1[910]^L1[905], L1[909]^L1[904]^L1[907], L1[908]^L1[907] };
	assign out[451:448]   = { L1[899]^L1[902]^L1[897], L1[898]^L1[901]^L1[896]^L1[899], L1[897]^L1[900]^L1[899]^L1[903]^L1[898], L1[896]^L1[903]^L1[898] };
	assign out[447:444]   = { L1[895]^L1[890], L1[894]^L1[889], L1[893]^L1[888]^L1[891], L1[892]^L1[891] };
	assign out[443:440]   = { L1[883]^L1[886]^L1[881], L1[882]^L1[885]^L1[880]^L1[883], L1[881]^L1[884]^L1[883]^L1[887]^L1[882], L1[880]^L1[887]^L1[882] };
	assign out[439:436]   = { L1[879]^L1[874], L1[878]^L1[873], L1[877]^L1[872]^L1[875], L1[876]^L1[875] };
	assign out[435:432]   = { L1[867]^L1[870]^L1[865], L1[866]^L1[869]^L1[864]^L1[867], L1[865]^L1[868]^L1[867]^L1[871]^L1[866], L1[864]^L1[871]^L1[866] };
	assign out[431:428]   = { L1[863]^L1[858], L1[862]^L1[857], L1[861]^L1[856]^L1[859], L1[860]^L1[859] };
	assign out[427:424]   = { L1[851]^L1[854]^L1[849], L1[850]^L1[853]^L1[848]^L1[851], L1[849]^L1[852]^L1[851]^L1[855]^L1[850], L1[848]^L1[855]^L1[850] };
	assign out[423:420]   = { L1[847]^L1[842], L1[846]^L1[841], L1[845]^L1[840]^L1[843], L1[844]^L1[843] };
	assign out[419:416]   = { L1[835]^L1[838]^L1[833], L1[834]^L1[837]^L1[832]^L1[835], L1[833]^L1[836]^L1[835]^L1[839]^L1[834], L1[832]^L1[839]^L1[834] };
	assign out[415:412]   = { L1[831]^L1[826], L1[830]^L1[825], L1[829]^L1[824]^L1[827], L1[828]^L1[827] };
	assign out[411:408]   = { L1[819]^L1[822]^L1[817], L1[818]^L1[821]^L1[816]^L1[819], L1[817]^L1[820]^L1[819]^L1[823]^L1[818], L1[816]^L1[823]^L1[818] };
	assign out[407:404]   = { L1[815]^L1[810], L1[814]^L1[809], L1[813]^L1[808]^L1[811], L1[812]^L1[811] };
	assign out[403:400]   = { L1[803]^L1[806]^L1[801], L1[802]^L1[805]^L1[800]^L1[803], L1[801]^L1[804]^L1[803]^L1[807]^L1[802], L1[800]^L1[807]^L1[802] };
	assign out[399:396]   = { L1[799]^L1[794], L1[798]^L1[793], L1[797]^L1[792]^L1[795], L1[796]^L1[795] };
	assign out[395:392]   = { L1[787]^L1[790]^L1[785], L1[786]^L1[789]^L1[784]^L1[787], L1[785]^L1[788]^L1[787]^L1[791]^L1[786], L1[784]^L1[791]^L1[786] };
	assign out[391:388]   = { L1[783]^L1[778], L1[782]^L1[777], L1[781]^L1[776]^L1[779], L1[780]^L1[779] };
	assign out[387:384]   = { L1[771]^L1[774]^L1[769], L1[770]^L1[773]^L1[768]^L1[771], L1[769]^L1[772]^L1[771]^L1[775]^L1[770], L1[768]^L1[775]^L1[770] };
	assign out[383:380]   = { L1[767]^L1[762], L1[766]^L1[761], L1[765]^L1[760]^L1[763], L1[764]^L1[763] };
	assign out[379:376]   = { L1[755]^L1[758]^L1[753], L1[754]^L1[757]^L1[752]^L1[755], L1[753]^L1[756]^L1[755]^L1[759]^L1[754], L1[752]^L1[759]^L1[754] };
	assign out[375:372]   = { L1[751]^L1[746], L1[750]^L1[745], L1[749]^L1[744]^L1[747], L1[748]^L1[747] };
	assign out[371:368]   = { L1[739]^L1[742]^L1[737], L1[738]^L1[741]^L1[736]^L1[739], L1[737]^L1[740]^L1[739]^L1[743]^L1[738], L1[736]^L1[743]^L1[738] };
	assign out[367:364]   = { L1[735]^L1[730], L1[734]^L1[729], L1[733]^L1[728]^L1[731], L1[732]^L1[731] };
	assign out[363:360]   = { L1[723]^L1[726]^L1[721], L1[722]^L1[725]^L1[720]^L1[723], L1[721]^L1[724]^L1[723]^L1[727]^L1[722], L1[720]^L1[727]^L1[722] };
	assign out[359:356]   = { L1[719]^L1[714], L1[718]^L1[713], L1[717]^L1[712]^L1[715], L1[716]^L1[715] };
	assign out[355:352]   = { L1[707]^L1[710]^L1[705], L1[706]^L1[709]^L1[704]^L1[707], L1[705]^L1[708]^L1[707]^L1[711]^L1[706], L1[704]^L1[711]^L1[706] };
	assign out[351:348]   = { L1[703]^L1[698], L1[702]^L1[697], L1[701]^L1[696]^L1[699], L1[700]^L1[699] };
	assign out[347:344]   = { L1[691]^L1[694]^L1[689], L1[690]^L1[693]^L1[688]^L1[691], L1[689]^L1[692]^L1[691]^L1[695]^L1[690], L1[688]^L1[695]^L1[690] };
	assign out[343:340]   = { L1[687]^L1[682], L1[686]^L1[681], L1[685]^L1[680]^L1[683], L1[684]^L1[683] };
	assign out[339:336]   = { L1[675]^L1[678]^L1[673], L1[674]^L1[677]^L1[672]^L1[675], L1[673]^L1[676]^L1[675]^L1[679]^L1[674], L1[672]^L1[679]^L1[674] };
	assign out[335:332]   = { L1[671]^L1[666], L1[670]^L1[665], L1[669]^L1[664]^L1[667], L1[668]^L1[667] };
	assign out[331:328]   = { L1[659]^L1[662]^L1[657], L1[658]^L1[661]^L1[656]^L1[659], L1[657]^L1[660]^L1[659]^L1[663]^L1[658], L1[656]^L1[663]^L1[658] };
	assign out[327:324]   = { L1[655]^L1[650], L1[654]^L1[649], L1[653]^L1[648]^L1[651], L1[652]^L1[651] };
	assign out[323:320]   = { L1[643]^L1[646]^L1[641], L1[642]^L1[645]^L1[640]^L1[643], L1[641]^L1[644]^L1[643]^L1[647]^L1[642], L1[640]^L1[647]^L1[642] };
	assign out[319:316]   = { L1[639]^L1[634], L1[638]^L1[633], L1[637]^L1[632]^L1[635], L1[636]^L1[635] };
	assign out[315:312]   = { L1[627]^L1[630]^L1[625], L1[626]^L1[629]^L1[624]^L1[627], L1[625]^L1[628]^L1[627]^L1[631]^L1[626], L1[624]^L1[631]^L1[626] };
	assign out[311:308]   = { L1[623]^L1[618], L1[622]^L1[617], L1[621]^L1[616]^L1[619], L1[620]^L1[619] };
	assign out[307:304]   = { L1[611]^L1[614]^L1[609], L1[610]^L1[613]^L1[608]^L1[611], L1[609]^L1[612]^L1[611]^L1[615]^L1[610], L1[608]^L1[615]^L1[610] };
	assign out[303:300]   = { L1[607]^L1[602], L1[606]^L1[601], L1[605]^L1[600]^L1[603], L1[604]^L1[603] };
	assign out[299:296]   = { L1[595]^L1[598]^L1[593], L1[594]^L1[597]^L1[592]^L1[595], L1[593]^L1[596]^L1[595]^L1[599]^L1[594], L1[592]^L1[599]^L1[594] };
	assign out[295:292]   = { L1[591]^L1[586], L1[590]^L1[585], L1[589]^L1[584]^L1[587], L1[588]^L1[587] };
	assign out[291:288]   = { L1[579]^L1[582]^L1[577], L1[578]^L1[581]^L1[576]^L1[579], L1[577]^L1[580]^L1[579]^L1[583]^L1[578], L1[576]^L1[583]^L1[578] };
	assign out[287:284]   = { L1[575]^L1[570], L1[574]^L1[569], L1[573]^L1[568]^L1[571], L1[572]^L1[571] };
	assign out[283:280]   = { L1[563]^L1[566]^L1[561], L1[562]^L1[565]^L1[560]^L1[563], L1[561]^L1[564]^L1[563]^L1[567]^L1[562], L1[560]^L1[567]^L1[562] };
	assign out[279:276]   = { L1[559]^L1[554], L1[558]^L1[553], L1[557]^L1[552]^L1[555], L1[556]^L1[555] };
	assign out[275:272]   = { L1[547]^L1[550]^L1[545], L1[546]^L1[549]^L1[544]^L1[547], L1[545]^L1[548]^L1[547]^L1[551]^L1[546], L1[544]^L1[551]^L1[546] };
	assign out[271:268]   = { L1[543]^L1[538], L1[542]^L1[537], L1[541]^L1[536]^L1[539], L1[540]^L1[539] };
	assign out[267:264]   = { L1[531]^L1[534]^L1[529], L1[530]^L1[533]^L1[528]^L1[531], L1[529]^L1[532]^L1[531]^L1[535]^L1[530], L1[528]^L1[535]^L1[530] };
	assign out[263:260]   = { L1[527]^L1[522], L1[526]^L1[521], L1[525]^L1[520]^L1[523], L1[524]^L1[523] };
	assign out[259:256]   = { L1[515]^L1[518]^L1[513], L1[514]^L1[517]^L1[512]^L1[515], L1[513]^L1[516]^L1[515]^L1[519]^L1[514], L1[512]^L1[519]^L1[514] };
	assign out[255:252]   = { L1[511]^L1[506], L1[510]^L1[505], L1[509]^L1[504]^L1[507], L1[508]^L1[507] };
	assign out[251:248]   = { L1[499]^L1[502]^L1[497], L1[498]^L1[501]^L1[496]^L1[499], L1[497]^L1[500]^L1[499]^L1[503]^L1[498], L1[496]^L1[503]^L1[498] };
	assign out[247:244]   = { L1[495]^L1[490], L1[494]^L1[489], L1[493]^L1[488]^L1[491], L1[492]^L1[491] };
	assign out[243:240]   = { L1[483]^L1[486]^L1[481], L1[482]^L1[485]^L1[480]^L1[483], L1[481]^L1[484]^L1[483]^L1[487]^L1[482], L1[480]^L1[487]^L1[482] };
	assign out[239:236]   = { L1[479]^L1[474], L1[478]^L1[473], L1[477]^L1[472]^L1[475], L1[476]^L1[475] };
	assign out[235:232]   = { L1[467]^L1[470]^L1[465], L1[466]^L1[469]^L1[464]^L1[467], L1[465]^L1[468]^L1[467]^L1[471]^L1[466], L1[464]^L1[471]^L1[466] };
	assign out[231:228]   = { L1[463]^L1[458], L1[462]^L1[457], L1[461]^L1[456]^L1[459], L1[460]^L1[459] };
	assign out[227:224]   = { L1[451]^L1[454]^L1[449], L1[450]^L1[453]^L1[448]^L1[451], L1[449]^L1[452]^L1[451]^L1[455]^L1[450], L1[448]^L1[455]^L1[450] };
	assign out[223:220]   = { L1[447]^L1[442], L1[446]^L1[441], L1[445]^L1[440]^L1[443], L1[444]^L1[443] };
	assign out[219:216]   = { L1[435]^L1[438]^L1[433], L1[434]^L1[437]^L1[432]^L1[435], L1[433]^L1[436]^L1[435]^L1[439]^L1[434], L1[432]^L1[439]^L1[434] };
	assign out[215:212]   = { L1[431]^L1[426], L1[430]^L1[425], L1[429]^L1[424]^L1[427], L1[428]^L1[427] };
	assign out[211:208]   = { L1[419]^L1[422]^L1[417], L1[418]^L1[421]^L1[416]^L1[419], L1[417]^L1[420]^L1[419]^L1[423]^L1[418], L1[416]^L1[423]^L1[418] };
	assign out[207:204]   = { L1[415]^L1[410], L1[414]^L1[409], L1[413]^L1[408]^L1[411], L1[412]^L1[411] };
	assign out[203:200]   = { L1[403]^L1[406]^L1[401], L1[402]^L1[405]^L1[400]^L1[403], L1[401]^L1[404]^L1[403]^L1[407]^L1[402], L1[400]^L1[407]^L1[402] };
	assign out[199:196]   = { L1[399]^L1[394], L1[398]^L1[393], L1[397]^L1[392]^L1[395], L1[396]^L1[395] };
	assign out[195:192]   = { L1[387]^L1[390]^L1[385], L1[386]^L1[389]^L1[384]^L1[387], L1[385]^L1[388]^L1[387]^L1[391]^L1[386], L1[384]^L1[391]^L1[386] };
	assign out[191:188]   = { L1[383]^L1[378], L1[382]^L1[377], L1[381]^L1[376]^L1[379], L1[380]^L1[379] };
	assign out[187:184]   = { L1[371]^L1[374]^L1[369], L1[370]^L1[373]^L1[368]^L1[371], L1[369]^L1[372]^L1[371]^L1[375]^L1[370], L1[368]^L1[375]^L1[370] };
	assign out[183:180]   = { L1[367]^L1[362], L1[366]^L1[361], L1[365]^L1[360]^L1[363], L1[364]^L1[363] };
	assign out[179:176]   = { L1[355]^L1[358]^L1[353], L1[354]^L1[357]^L1[352]^L1[355], L1[353]^L1[356]^L1[355]^L1[359]^L1[354], L1[352]^L1[359]^L1[354] };
	assign out[175:172]   = { L1[351]^L1[346], L1[350]^L1[345], L1[349]^L1[344]^L1[347], L1[348]^L1[347] };
	assign out[171:168]   = { L1[339]^L1[342]^L1[337], L1[338]^L1[341]^L1[336]^L1[339], L1[337]^L1[340]^L1[339]^L1[343]^L1[338], L1[336]^L1[343]^L1[338] };
	assign out[167:164]   = { L1[335]^L1[330], L1[334]^L1[329], L1[333]^L1[328]^L1[331], L1[332]^L1[331] };
	assign out[163:160]   = { L1[323]^L1[326]^L1[321], L1[322]^L1[325]^L1[320]^L1[323], L1[321]^L1[324]^L1[323]^L1[327]^L1[322], L1[320]^L1[327]^L1[322] };
	assign out[159:156]   = { L1[319]^L1[314], L1[318]^L1[313], L1[317]^L1[312]^L1[315], L1[316]^L1[315] };
	assign out[155:152]   = { L1[307]^L1[310]^L1[305], L1[306]^L1[309]^L1[304]^L1[307], L1[305]^L1[308]^L1[307]^L1[311]^L1[306], L1[304]^L1[311]^L1[306] };
	assign out[151:148]   = { L1[303]^L1[298], L1[302]^L1[297], L1[301]^L1[296]^L1[299], L1[300]^L1[299] };
	assign out[147:144]   = { L1[291]^L1[294]^L1[289], L1[290]^L1[293]^L1[288]^L1[291], L1[289]^L1[292]^L1[291]^L1[295]^L1[290], L1[288]^L1[295]^L1[290] };
	assign out[143:140]   = { L1[287]^L1[282], L1[286]^L1[281], L1[285]^L1[280]^L1[283], L1[284]^L1[283] };
	assign out[139:136]   = { L1[275]^L1[278]^L1[273], L1[274]^L1[277]^L1[272]^L1[275], L1[273]^L1[276]^L1[275]^L1[279]^L1[274], L1[272]^L1[279]^L1[274] };
	assign out[135:132]   = { L1[271]^L1[266], L1[270]^L1[265], L1[269]^L1[264]^L1[267], L1[268]^L1[267] };
	assign out[131:128]   = { L1[259]^L1[262]^L1[257], L1[258]^L1[261]^L1[256]^L1[259], L1[257]^L1[260]^L1[259]^L1[263]^L1[258], L1[256]^L1[263]^L1[258] };
	assign out[127:124]   = { L1[255]^L1[250], L1[254]^L1[249], L1[253]^L1[248]^L1[251], L1[252]^L1[251] };
	assign out[123:120]   = { L1[243]^L1[246]^L1[241], L1[242]^L1[245]^L1[240]^L1[243], L1[241]^L1[244]^L1[243]^L1[247]^L1[242], L1[240]^L1[247]^L1[242] };
	assign out[119:116]   = { L1[239]^L1[234], L1[238]^L1[233], L1[237]^L1[232]^L1[235], L1[236]^L1[235] };
	assign out[115:112]   = { L1[227]^L1[230]^L1[225], L1[226]^L1[229]^L1[224]^L1[227], L1[225]^L1[228]^L1[227]^L1[231]^L1[226], L1[224]^L1[231]^L1[226] };
	assign out[111:108]   = { L1[223]^L1[218], L1[222]^L1[217], L1[221]^L1[216]^L1[219], L1[220]^L1[219] };
	assign out[107:104]   = { L1[211]^L1[214]^L1[209], L1[210]^L1[213]^L1[208]^L1[211], L1[209]^L1[212]^L1[211]^L1[215]^L1[210], L1[208]^L1[215]^L1[210] };
	assign out[103:100]   = { L1[207]^L1[202], L1[206]^L1[201], L1[205]^L1[200]^L1[203], L1[204]^L1[203] };
	assign out[ 99: 96]   = { L1[195]^L1[198]^L1[193], L1[194]^L1[197]^L1[192]^L1[195], L1[193]^L1[196]^L1[195]^L1[199]^L1[194], L1[192]^L1[199]^L1[194] };
	assign out[ 95: 92]   = { L1[191]^L1[186], L1[190]^L1[185], L1[189]^L1[184]^L1[187], L1[188]^L1[187] };
	assign out[ 91: 88]   = { L1[179]^L1[182]^L1[177], L1[178]^L1[181]^L1[176]^L1[179], L1[177]^L1[180]^L1[179]^L1[183]^L1[178], L1[176]^L1[183]^L1[178] };
	assign out[ 87: 84]   = { L1[175]^L1[170], L1[174]^L1[169], L1[173]^L1[168]^L1[171], L1[172]^L1[171] };
	assign out[ 83: 80]   = { L1[163]^L1[166]^L1[161], L1[162]^L1[165]^L1[160]^L1[163], L1[161]^L1[164]^L1[163]^L1[167]^L1[162], L1[160]^L1[167]^L1[162] };
	assign out[ 79: 76]   = { L1[159]^L1[154], L1[158]^L1[153], L1[157]^L1[152]^L1[155], L1[156]^L1[155] };
	assign out[ 75: 72]   = { L1[147]^L1[150]^L1[145], L1[146]^L1[149]^L1[144]^L1[147], L1[145]^L1[148]^L1[147]^L1[151]^L1[146], L1[144]^L1[151]^L1[146] };
	assign out[ 71: 68]   = { L1[143]^L1[138], L1[142]^L1[137], L1[141]^L1[136]^L1[139], L1[140]^L1[139] };
	assign out[ 67: 64]   = { L1[131]^L1[134]^L1[129], L1[130]^L1[133]^L1[128]^L1[131], L1[129]^L1[132]^L1[131]^L1[135]^L1[130], L1[128]^L1[135]^L1[130] };
	assign out[ 63: 60]   = { L1[127]^L1[122], L1[126]^L1[121], L1[125]^L1[120]^L1[123], L1[124]^L1[123] };
	assign out[ 59: 56]   = { L1[115]^L1[118]^L1[113], L1[114]^L1[117]^L1[112]^L1[115], L1[113]^L1[116]^L1[115]^L1[119]^L1[114], L1[112]^L1[119]^L1[114] };
	assign out[ 55: 52]   = { L1[111]^L1[106], L1[110]^L1[105], L1[109]^L1[104]^L1[107], L1[108]^L1[107] };
	assign out[ 51: 48]   = { L1[99]^L1[102]^L1[97], L1[98]^L1[101]^L1[96]^L1[99], L1[97]^L1[100]^L1[99]^L1[103]^L1[98], L1[96]^L1[103]^L1[98] };
	assign out[ 47: 44]   = { L1[95]^L1[90], L1[94]^L1[89], L1[93]^L1[88]^L1[91], L1[92]^L1[91] };
	assign out[ 43: 40]   = { L1[83]^L1[86]^L1[81], L1[82]^L1[85]^L1[80]^L1[83], L1[81]^L1[84]^L1[83]^L1[87]^L1[82], L1[80]^L1[87]^L1[82] };
	assign out[ 39: 36]   = { L1[79]^L1[74], L1[78]^L1[73], L1[77]^L1[72]^L1[75], L1[76]^L1[75] };
	assign out[ 35: 32]   = { L1[67]^L1[70]^L1[65], L1[66]^L1[69]^L1[64]^L1[67], L1[65]^L1[68]^L1[67]^L1[71]^L1[66], L1[64]^L1[71]^L1[66] };
	assign out[ 31: 28]   = { L1[63]^L1[58], L1[62]^L1[57], L1[61]^L1[56]^L1[59], L1[60]^L1[59] };
	assign out[ 27: 24]   = { L1[51]^L1[54]^L1[49], L1[50]^L1[53]^L1[48]^L1[51], L1[49]^L1[52]^L1[51]^L1[55]^L1[50], L1[48]^L1[55]^L1[50] };
	assign out[ 23: 20]   = { L1[47]^L1[42], L1[46]^L1[41], L1[45]^L1[40]^L1[43], L1[44]^L1[43] };
	assign out[ 19: 16]   = { L1[35]^L1[38]^L1[33], L1[34]^L1[37]^L1[32]^L1[35], L1[33]^L1[36]^L1[35]^L1[39]^L1[34], L1[32]^L1[39]^L1[34] };
	assign out[ 15: 12]   = { L1[31]^L1[26], L1[30]^L1[25], L1[29]^L1[24]^L1[27], L1[28]^L1[27] };
	assign out[ 11:  8]   = { L1[19]^L1[22]^L1[17], L1[18]^L1[21]^L1[16]^L1[19], L1[17]^L1[20]^L1[19]^L1[23]^L1[18], L1[16]^L1[23]^L1[18] };
	assign out[  7:  4]   = { L1[15]^L1[10], L1[14]^L1[9], L1[13]^L1[8]^L1[11], L1[12]^L1[11] };
	assign out[  3:  0]   = { L1[3]^L1[6]^L1[1], L1[2]^L1[5]^L1[0]^L1[3], L1[1]^L1[4]^L1[3]^L1[7]^L1[2], L1[0]^L1[7]^L1[2] };

endmodule 

module jh_round_b (
	input [255:0] in, 
	output [255:0] out
);

	wire [3:0] sbox [0:15] = { 4'h9,4'h1,4'hd,4'h7,4'h4,4'h2,4'h3,4'h8,4'h0,4'ha,4'hc,4'h5,4'hb,4'h6,4'hf,4'he };

	wire [255:0] L1;

	assign L1[255:252] = sbox[ in[255:252] ];
	assign L1[251:248] = sbox[ in[251:248] ];
	assign L1[247:244] = sbox[ in[247:244] ];
	assign L1[243:240] = sbox[ in[243:240] ];
	assign L1[239:236] = sbox[ in[239:236] ];
	assign L1[235:232] = sbox[ in[235:232] ];
	assign L1[231:228] = sbox[ in[231:228] ];
	assign L1[227:224] = sbox[ in[227:224] ];
	assign L1[223:220] = sbox[ in[223:220] ];
	assign L1[219:216] = sbox[ in[219:216] ];
	assign L1[215:212] = sbox[ in[215:212] ];
	assign L1[211:208] = sbox[ in[211:208] ];
	assign L1[207:204] = sbox[ in[207:204] ];
	assign L1[203:200] = sbox[ in[203:200] ];
	assign L1[199:196] = sbox[ in[199:196] ];
	assign L1[195:192] = sbox[ in[195:192] ];
	assign L1[191:188] = sbox[ in[191:188] ];
	assign L1[187:184] = sbox[ in[187:184] ];
	assign L1[183:180] = sbox[ in[183:180] ];
	assign L1[179:176] = sbox[ in[179:176] ];
	assign L1[175:172] = sbox[ in[175:172] ];
	assign L1[171:168] = sbox[ in[171:168] ];
	assign L1[167:164] = sbox[ in[167:164] ];
	assign L1[163:160] = sbox[ in[163:160] ];
	assign L1[159:156] = sbox[ in[159:156] ];
	assign L1[155:152] = sbox[ in[155:152] ];
	assign L1[151:148] = sbox[ in[151:148] ];
	assign L1[147:144] = sbox[ in[147:144] ];
	assign L1[143:140] = sbox[ in[143:140] ];
	assign L1[139:136] = sbox[ in[139:136] ];
	assign L1[135:132] = sbox[ in[135:132] ];
	assign L1[131:128] = sbox[ in[131:128] ];
	assign L1[127:124] = sbox[ in[127:124] ];
	assign L1[123:120] = sbox[ in[123:120] ];
	assign L1[119:116] = sbox[ in[119:116] ];
	assign L1[115:112] = sbox[ in[115:112] ];
	assign L1[111:108] = sbox[ in[111:108] ];
	assign L1[107:104] = sbox[ in[107:104] ];
	assign L1[103:100] = sbox[ in[103:100] ];
	assign L1[99:96] = sbox[ in[99:96] ];
	assign L1[95:92] = sbox[ in[95:92] ];
	assign L1[91:88] = sbox[ in[91:88] ];
	assign L1[87:84] = sbox[ in[87:84] ];
	assign L1[83:80] = sbox[ in[83:80] ];
	assign L1[79:76] = sbox[ in[79:76] ];
	assign L1[75:72] = sbox[ in[75:72] ];
	assign L1[71:68] = sbox[ in[71:68] ];
	assign L1[67:64] = sbox[ in[67:64] ];
	assign L1[63:60] = sbox[ in[63:60] ];
	assign L1[59:56] = sbox[ in[59:56] ];
	assign L1[55:52] = sbox[ in[55:52] ];
	assign L1[51:48] = sbox[ in[51:48] ];
	assign L1[47:44] = sbox[ in[47:44] ];
	assign L1[43:40] = sbox[ in[43:40] ];
	assign L1[39:36] = sbox[ in[39:36] ];
	assign L1[35:32] = sbox[ in[35:32] ];
	assign L1[31:28] = sbox[ in[31:28] ];
	assign L1[27:24] = sbox[ in[27:24] ];
	assign L1[23:20] = sbox[ in[23:20] ];
	assign L1[19:16] = sbox[ in[19:16] ];
	assign L1[15:12] = sbox[ in[15:12] ];
	assign L1[11:8] = sbox[ in[11:8] ];
	assign L1[7:4] = sbox[ in[7:4] ];
	assign L1[3:0] = sbox[ in[3:0] ];

	assign out[255:252] = { L1[244]^L1[243], L1[245]^L1[240]^L1[243], L1[246]^L1[241], L1[247]^L1[242] };
	assign out[251:248] = { L1[248]^L1[255]^L1[250], L1[249]^L1[252]^L1[251]^L1[255]^L1[250], L1[250]^L1[253]^L1[248]^L1[251], L1[251]^L1[254]^L1[249] };
	assign out[247:244] = { L1[228]^L1[227], L1[229]^L1[224]^L1[227], L1[230]^L1[225], L1[231]^L1[226] };
	assign out[243:240] = { L1[232]^L1[239]^L1[234], L1[233]^L1[236]^L1[235]^L1[239]^L1[234], L1[234]^L1[237]^L1[232]^L1[235], L1[235]^L1[238]^L1[233] };
	assign out[239:236] = { L1[212]^L1[211], L1[213]^L1[208]^L1[211], L1[214]^L1[209], L1[215]^L1[210] };
	assign out[235:232] = { L1[216]^L1[223]^L1[218], L1[217]^L1[220]^L1[219]^L1[223]^L1[218], L1[218]^L1[221]^L1[216]^L1[219], L1[219]^L1[222]^L1[217] };
	assign out[231:228] = { L1[196]^L1[195], L1[197]^L1[192]^L1[195], L1[198]^L1[193], L1[199]^L1[194] };
	assign out[227:224] = { L1[200]^L1[207]^L1[202], L1[201]^L1[204]^L1[203]^L1[207]^L1[202], L1[202]^L1[205]^L1[200]^L1[203], L1[203]^L1[206]^L1[201] };
	assign out[223:220] = { L1[180]^L1[179], L1[181]^L1[176]^L1[179], L1[182]^L1[177], L1[183]^L1[178] };
	assign out[219:216] = { L1[184]^L1[191]^L1[186], L1[185]^L1[188]^L1[187]^L1[191]^L1[186], L1[186]^L1[189]^L1[184]^L1[187], L1[187]^L1[190]^L1[185] };
	assign out[215:212] = { L1[164]^L1[163], L1[165]^L1[160]^L1[163], L1[166]^L1[161], L1[167]^L1[162] };
	assign out[211:208] = { L1[168]^L1[175]^L1[170], L1[169]^L1[172]^L1[171]^L1[175]^L1[170], L1[170]^L1[173]^L1[168]^L1[171], L1[171]^L1[174]^L1[169] };
	assign out[207:204] = { L1[148]^L1[147], L1[149]^L1[144]^L1[147], L1[150]^L1[145], L1[151]^L1[146] };
	assign out[203:200] = { L1[152]^L1[159]^L1[154], L1[153]^L1[156]^L1[155]^L1[159]^L1[154], L1[154]^L1[157]^L1[152]^L1[155], L1[155]^L1[158]^L1[153] };
	assign out[199:196] = { L1[132]^L1[131], L1[133]^L1[128]^L1[131], L1[134]^L1[129], L1[135]^L1[130] };
	assign out[195:192] = { L1[136]^L1[143]^L1[138], L1[137]^L1[140]^L1[139]^L1[143]^L1[138], L1[138]^L1[141]^L1[136]^L1[139], L1[139]^L1[142]^L1[137] };
	assign out[191:188] = { L1[116]^L1[115], L1[117]^L1[112]^L1[115], L1[118]^L1[113], L1[119]^L1[114] };
	assign out[187:184] = { L1[120]^L1[127]^L1[122], L1[121]^L1[124]^L1[123]^L1[127]^L1[122], L1[122]^L1[125]^L1[120]^L1[123], L1[123]^L1[126]^L1[121] };
	assign out[183:180] = { L1[100]^L1[99], L1[101]^L1[96]^L1[99], L1[102]^L1[97], L1[103]^L1[98] };
	assign out[179:176] = { L1[104]^L1[111]^L1[106], L1[105]^L1[108]^L1[107]^L1[111]^L1[106], L1[106]^L1[109]^L1[104]^L1[107], L1[107]^L1[110]^L1[105] };
	assign out[175:172] = { L1[84]^L1[83], L1[85]^L1[80]^L1[83], L1[86]^L1[81], L1[87]^L1[82] };
	assign out[171:168] = { L1[88]^L1[95]^L1[90], L1[89]^L1[92]^L1[91]^L1[95]^L1[90], L1[90]^L1[93]^L1[88]^L1[91], L1[91]^L1[94]^L1[89] };
	assign out[167:164] = { L1[68]^L1[67], L1[69]^L1[64]^L1[67], L1[70]^L1[65], L1[71]^L1[66] };
	assign out[163:160] = { L1[72]^L1[79]^L1[74], L1[73]^L1[76]^L1[75]^L1[79]^L1[74], L1[74]^L1[77]^L1[72]^L1[75], L1[75]^L1[78]^L1[73] };
	assign out[159:156] = { L1[52]^L1[51], L1[53]^L1[48]^L1[51], L1[54]^L1[49], L1[55]^L1[50] };
	assign out[155:152] = { L1[56]^L1[63]^L1[58], L1[57]^L1[60]^L1[59]^L1[63]^L1[58], L1[58]^L1[61]^L1[56]^L1[59], L1[59]^L1[62]^L1[57] };
	assign out[151:148] = { L1[36]^L1[35], L1[37]^L1[32]^L1[35], L1[38]^L1[33], L1[39]^L1[34] };
	assign out[147:144] = { L1[40]^L1[47]^L1[42], L1[41]^L1[44]^L1[43]^L1[47]^L1[42], L1[42]^L1[45]^L1[40]^L1[43], L1[43]^L1[46]^L1[41] };
	assign out[143:140] = { L1[20]^L1[19], L1[21]^L1[16]^L1[19], L1[22]^L1[17], L1[23]^L1[18] };
	assign out[139:136] = { L1[24]^L1[31]^L1[26], L1[25]^L1[28]^L1[27]^L1[31]^L1[26], L1[26]^L1[29]^L1[24]^L1[27], L1[27]^L1[30]^L1[25] };
	assign out[135:132] = { L1[4]^L1[3], L1[5]^L1[0]^L1[3], L1[6]^L1[1], L1[7]^L1[2] };
	assign out[131:128] = { L1[8]^L1[15]^L1[10], L1[9]^L1[12]^L1[11]^L1[15]^L1[10], L1[10]^L1[13]^L1[8]^L1[11], L1[11]^L1[14]^L1[9] };
	assign out[127:124] = { L1[252]^L1[251], L1[253]^L1[248]^L1[251], L1[254]^L1[249], L1[255]^L1[250] };
	assign out[123:120] = { L1[240]^L1[247]^L1[242], L1[241]^L1[244]^L1[243]^L1[247]^L1[242], L1[242]^L1[245]^L1[240]^L1[243], L1[243]^L1[246]^L1[241] };
	assign out[119:116] = { L1[236]^L1[235], L1[237]^L1[232]^L1[235], L1[238]^L1[233], L1[239]^L1[234] };
	assign out[115:112] = { L1[224]^L1[231]^L1[226], L1[225]^L1[228]^L1[227]^L1[231]^L1[226], L1[226]^L1[229]^L1[224]^L1[227], L1[227]^L1[230]^L1[225] };
	assign out[111:108] = { L1[220]^L1[219], L1[221]^L1[216]^L1[219], L1[222]^L1[217], L1[223]^L1[218] };
	assign out[107:104] = { L1[208]^L1[215]^L1[210], L1[209]^L1[212]^L1[211]^L1[215]^L1[210], L1[210]^L1[213]^L1[208]^L1[211], L1[211]^L1[214]^L1[209] };
	assign out[103:100] = { L1[204]^L1[203], L1[205]^L1[200]^L1[203], L1[206]^L1[201], L1[207]^L1[202] };
	assign out[99:96]   = { L1[192]^L1[199]^L1[194], L1[193]^L1[196]^L1[195]^L1[199]^L1[194], L1[194]^L1[197]^L1[192]^L1[195], L1[195]^L1[198]^L1[193] };
	assign out[95:92]   = { L1[188]^L1[187], L1[189]^L1[184]^L1[187], L1[190]^L1[185], L1[191]^L1[186] };
	assign out[91:88]   = { L1[176]^L1[183]^L1[178], L1[177]^L1[180]^L1[179]^L1[183]^L1[178], L1[178]^L1[181]^L1[176]^L1[179], L1[179]^L1[182]^L1[177] };
	assign out[87:84]   = { L1[172]^L1[171], L1[173]^L1[168]^L1[171], L1[174]^L1[169], L1[175]^L1[170] };
	assign out[83:80]   = { L1[160]^L1[167]^L1[162], L1[161]^L1[164]^L1[163]^L1[167]^L1[162], L1[162]^L1[165]^L1[160]^L1[163], L1[163]^L1[166]^L1[161] };
	assign out[79:76]   = { L1[156]^L1[155], L1[157]^L1[152]^L1[155], L1[158]^L1[153], L1[159]^L1[154] };
	assign out[75:72]   = { L1[144]^L1[151]^L1[146], L1[145]^L1[148]^L1[147]^L1[151]^L1[146], L1[146]^L1[149]^L1[144]^L1[147], L1[147]^L1[150]^L1[145] };
	assign out[71:68]   = { L1[140]^L1[139], L1[141]^L1[136]^L1[139], L1[142]^L1[137], L1[143]^L1[138] };
	assign out[67:64]   = { L1[128]^L1[135]^L1[130], L1[129]^L1[132]^L1[131]^L1[135]^L1[130], L1[130]^L1[133]^L1[128]^L1[131], L1[131]^L1[134]^L1[129] };
	assign out[63:60]   = { L1[124]^L1[123], L1[125]^L1[120]^L1[123], L1[126]^L1[121], L1[127]^L1[122] };
	assign out[59:56]   = { L1[112]^L1[119]^L1[114], L1[113]^L1[116]^L1[115]^L1[119]^L1[114], L1[114]^L1[117]^L1[112]^L1[115], L1[115]^L1[118]^L1[113] };
	assign out[55:52]   = { L1[108]^L1[107], L1[109]^L1[104]^L1[107], L1[110]^L1[105], L1[111]^L1[106] };
	assign out[51:48]   = { L1[96]^L1[103]^L1[98], L1[97]^L1[100]^L1[99]^L1[103]^L1[98], L1[98]^L1[101]^L1[96]^L1[99], L1[99]^L1[102]^L1[97] };
	assign out[47:44]   = { L1[92]^L1[91], L1[93]^L1[88]^L1[91], L1[94]^L1[89], L1[95]^L1[90] };
	assign out[43:40]   = { L1[80]^L1[87]^L1[82], L1[81]^L1[84]^L1[83]^L1[87]^L1[82], L1[82]^L1[85]^L1[80]^L1[83], L1[83]^L1[86]^L1[81] };
	assign out[39:36]   = { L1[76]^L1[75], L1[77]^L1[72]^L1[75], L1[78]^L1[73], L1[79]^L1[74] };
	assign out[35:32]   = { L1[64]^L1[71]^L1[66], L1[65]^L1[68]^L1[67]^L1[71]^L1[66], L1[66]^L1[69]^L1[64]^L1[67], L1[67]^L1[70]^L1[65] };
	assign out[31:28]   = { L1[60]^L1[59], L1[61]^L1[56]^L1[59], L1[62]^L1[57], L1[63]^L1[58] };
	assign out[27:24]   = { L1[48]^L1[55]^L1[50], L1[49]^L1[52]^L1[51]^L1[55]^L1[50], L1[50]^L1[53]^L1[48]^L1[51], L1[51]^L1[54]^L1[49] };
	assign out[23:20]   = { L1[44]^L1[43], L1[45]^L1[40]^L1[43], L1[46]^L1[41], L1[47]^L1[42] };
	assign out[19:16]   = { L1[32]^L1[39]^L1[34], L1[33]^L1[36]^L1[35]^L1[39]^L1[34], L1[34]^L1[37]^L1[32]^L1[35], L1[35]^L1[38]^L1[33] };
	assign out[15:12]   = { L1[28]^L1[27], L1[29]^L1[24]^L1[27], L1[30]^L1[25], L1[31]^L1[26] };
	assign out[11:8]    = { L1[16]^L1[23]^L1[18], L1[17]^L1[20]^L1[19]^L1[23]^L1[18], L1[18]^L1[21]^L1[16]^L1[19], L1[19]^L1[22]^L1[17] };
	assign out[7:4]     = { L1[12]^L1[11], L1[13]^L1[8]^L1[11], L1[14]^L1[9], L1[15]^L1[10] };
	assign out[3:0]     = { L1[0]^L1[7]^L1[2], L1[1]^L1[4]^L1[3]^L1[7]^L1[2], L1[2]^L1[5]^L1[0]^L1[3], L1[3]^L1[6]^L1[1] };

endmodule 

module jh_final (
	input [1023:0] in,
	output [1023:0] out
);

	 assign { out[7], out[263], out[519], out[775] } = in[3:0];
	 assign { out[6], out[262], out[518], out[774] } = in[11:8];
	 assign { out[5], out[261], out[517], out[773] } = in[19:16];
	 assign { out[4], out[260], out[516], out[772] } = in[27:24];
	 assign { out[3], out[259], out[515], out[771] } = in[35:32];
	 assign { out[2], out[258], out[514], out[770] } = in[43:40];
	 assign { out[1], out[257], out[513], out[769] } = in[51:48];
	 assign { out[0], out[256], out[512], out[768] } = in[59:56];
	 assign { out[15], out[271], out[527], out[783] } = in[67:64];
	 assign { out[14], out[270], out[526], out[782] } = in[75:72];
	 assign { out[13], out[269], out[525], out[781] } = in[83:80];
	 assign { out[12], out[268], out[524], out[780] } = in[91:88];
	 assign { out[11], out[267], out[523], out[779] } = in[99:96];
	 assign { out[10], out[266], out[522], out[778] } = in[107:104];
	 assign { out[9], out[265], out[521], out[777] } = in[115:112];
	 assign { out[8], out[264], out[520], out[776] } = in[123:120];
	 assign { out[23], out[279], out[535], out[791] } = in[131:128];
	 assign { out[22], out[278], out[534], out[790] } = in[139:136];
	 assign { out[21], out[277], out[533], out[789] } = in[147:144];
	 assign { out[20], out[276], out[532], out[788] } = in[155:152];
	 assign { out[19], out[275], out[531], out[787] } = in[163:160];
	 assign { out[18], out[274], out[530], out[786] } = in[171:168];
	 assign { out[17], out[273], out[529], out[785] } = in[179:176];
	 assign { out[16], out[272], out[528], out[784] } = in[187:184];
	 assign { out[31], out[287], out[543], out[799] } = in[195:192];
	 assign { out[30], out[286], out[542], out[798] } = in[203:200];
	 assign { out[29], out[285], out[541], out[797] } = in[211:208];
	 assign { out[28], out[284], out[540], out[796] } = in[219:216];
	 assign { out[27], out[283], out[539], out[795] } = in[227:224];
	 assign { out[26], out[282], out[538], out[794] } = in[235:232];
	 assign { out[25], out[281], out[537], out[793] } = in[243:240];
	 assign { out[24], out[280], out[536], out[792] } = in[251:248];
	 assign { out[39], out[295], out[551], out[807] } = in[259:256];
	 assign { out[38], out[294], out[550], out[806] } = in[267:264];
	 assign { out[37], out[293], out[549], out[805] } = in[275:272];
	 assign { out[36], out[292], out[548], out[804] } = in[283:280];
	 assign { out[35], out[291], out[547], out[803] } = in[291:288];
	 assign { out[34], out[290], out[546], out[802] } = in[299:296];
	 assign { out[33], out[289], out[545], out[801] } = in[307:304];
	 assign { out[32], out[288], out[544], out[800] } = in[315:312];
	 assign { out[47], out[303], out[559], out[815] } = in[323:320];
	 assign { out[46], out[302], out[558], out[814] } = in[331:328];
	 assign { out[45], out[301], out[557], out[813] } = in[339:336];
	 assign { out[44], out[300], out[556], out[812] } = in[347:344];
	 assign { out[43], out[299], out[555], out[811] } = in[355:352];
	 assign { out[42], out[298], out[554], out[810] } = in[363:360];
	 assign { out[41], out[297], out[553], out[809] } = in[371:368];
	 assign { out[40], out[296], out[552], out[808] } = in[379:376];
	 assign { out[55], out[311], out[567], out[823] } = in[387:384];
	 assign { out[54], out[310], out[566], out[822] } = in[395:392];
	 assign { out[53], out[309], out[565], out[821] } = in[403:400];
	 assign { out[52], out[308], out[564], out[820] } = in[411:408];
	 assign { out[51], out[307], out[563], out[819] } = in[419:416];
	 assign { out[50], out[306], out[562], out[818] } = in[427:424];
	 assign { out[49], out[305], out[561], out[817] } = in[435:432];
	 assign { out[48], out[304], out[560], out[816] } = in[443:440];
	 assign { out[63], out[319], out[575], out[831] } = in[451:448];
	 assign { out[62], out[318], out[574], out[830] } = in[459:456];
	 assign { out[61], out[317], out[573], out[829] } = in[467:464];
	 assign { out[60], out[316], out[572], out[828] } = in[475:472];
	 assign { out[59], out[315], out[571], out[827] } = in[483:480];
	 assign { out[58], out[314], out[570], out[826] } = in[491:488];
	 assign { out[57], out[313], out[569], out[825] } = in[499:496];
	 assign { out[56], out[312], out[568], out[824] } = in[507:504];
	 assign { out[71], out[327], out[583], out[839] } = in[515:512];
	 assign { out[70], out[326], out[582], out[838] } = in[523:520];
	 assign { out[69], out[325], out[581], out[837] } = in[531:528];
	 assign { out[68], out[324], out[580], out[836] } = in[539:536];
	 assign { out[67], out[323], out[579], out[835] } = in[547:544];
	 assign { out[66], out[322], out[578], out[834] } = in[555:552];
	 assign { out[65], out[321], out[577], out[833] } = in[563:560];
	 assign { out[64], out[320], out[576], out[832] } = in[571:568];
	 assign { out[79], out[335], out[591], out[847] } = in[579:576];
	 assign { out[78], out[334], out[590], out[846] } = in[587:584];
	 assign { out[77], out[333], out[589], out[845] } = in[595:592];
	 assign { out[76], out[332], out[588], out[844] } = in[603:600];
	 assign { out[75], out[331], out[587], out[843] } = in[611:608];
	 assign { out[74], out[330], out[586], out[842] } = in[619:616];
	 assign { out[73], out[329], out[585], out[841] } = in[627:624];
	 assign { out[72], out[328], out[584], out[840] } = in[635:632];
	 assign { out[87], out[343], out[599], out[855] } = in[643:640];
	 assign { out[86], out[342], out[598], out[854] } = in[651:648];
	 assign { out[85], out[341], out[597], out[853] } = in[659:656];
	 assign { out[84], out[340], out[596], out[852] } = in[667:664];
	 assign { out[83], out[339], out[595], out[851] } = in[675:672];
	 assign { out[82], out[338], out[594], out[850] } = in[683:680];
	 assign { out[81], out[337], out[593], out[849] } = in[691:688];
	 assign { out[80], out[336], out[592], out[848] } = in[699:696];
	 assign { out[95], out[351], out[607], out[863] } = in[707:704];
	 assign { out[94], out[350], out[606], out[862] } = in[715:712];
	 assign { out[93], out[349], out[605], out[861] } = in[723:720];
	 assign { out[92], out[348], out[604], out[860] } = in[731:728];
	 assign { out[91], out[347], out[603], out[859] } = in[739:736];
	 assign { out[90], out[346], out[602], out[858] } = in[747:744];
	 assign { out[89], out[345], out[601], out[857] } = in[755:752];
	 assign { out[88], out[344], out[600], out[856] } = in[763:760];
	 assign { out[103], out[359], out[615], out[871] } = in[771:768];
	 assign { out[102], out[358], out[614], out[870] } = in[779:776];
	 assign { out[101], out[357], out[613], out[869] } = in[787:784];
	 assign { out[100], out[356], out[612], out[868] } = in[795:792];
	 assign { out[99], out[355], out[611], out[867] } = in[803:800];
	 assign { out[98], out[354], out[610], out[866] } = in[811:808];
	 assign { out[97], out[353], out[609], out[865] } = in[819:816];
	 assign { out[96], out[352], out[608], out[864] } = in[827:824];
	 assign { out[111], out[367], out[623], out[879] } = in[835:832];
	 assign { out[110], out[366], out[622], out[878] } = in[843:840];
	 assign { out[109], out[365], out[621], out[877] } = in[851:848];
	 assign { out[108], out[364], out[620], out[876] } = in[859:856];
	 assign { out[107], out[363], out[619], out[875] } = in[867:864];
	 assign { out[106], out[362], out[618], out[874] } = in[875:872];
	 assign { out[105], out[361], out[617], out[873] } = in[883:880];
	 assign { out[104], out[360], out[616], out[872] } = in[891:888];
	 assign { out[119], out[375], out[631], out[887] } = in[899:896];
	 assign { out[118], out[374], out[630], out[886] } = in[907:904];
	 assign { out[117], out[373], out[629], out[885] } = in[915:912];
	 assign { out[116], out[372], out[628], out[884] } = in[923:920];
	 assign { out[115], out[371], out[627], out[883] } = in[931:928];
	 assign { out[114], out[370], out[626], out[882] } = in[939:936];
	 assign { out[113], out[369], out[625], out[881] } = in[947:944];
	 assign { out[112], out[368], out[624], out[880] } = in[955:952];
	 assign { out[127], out[383], out[639], out[895] } = in[963:960];
	 assign { out[126], out[382], out[638], out[894] } = in[971:968];
	 assign { out[125], out[381], out[637], out[893] } = in[979:976];
	 assign { out[124], out[380], out[636], out[892] } = in[987:984];
	 assign { out[123], out[379], out[635], out[891] } = in[995:992];
	 assign { out[122], out[378], out[634], out[890] } = in[1003:1000];
	 assign { out[121], out[377], out[633], out[889] } = in[1011:1008];
	 assign { out[120], out[376], out[632], out[888] } = in[1019:1016];
	 assign { out[135], out[391], out[647], out[903] } = in[7:4];
	 assign { out[134], out[390], out[646], out[902] } = in[15:12];
	 assign { out[133], out[389], out[645], out[901] } = in[23:20];
	 assign { out[132], out[388], out[644], out[900] } = in[31:28];
	 assign { out[131], out[387], out[643], out[899] } = in[39:36];
	 assign { out[130], out[386], out[642], out[898] } = in[47:44];
	 assign { out[129], out[385], out[641], out[897] } = in[55:52];
	 assign { out[128], out[384], out[640], out[896] } = in[63:60];
	 assign { out[143], out[399], out[655], out[911] } = in[71:68];
	 assign { out[142], out[398], out[654], out[910] } = in[79:76];
	 assign { out[141], out[397], out[653], out[909] } = in[87:84];
	 assign { out[140], out[396], out[652], out[908] } = in[95:92];
	 assign { out[139], out[395], out[651], out[907] } = in[103:100];
	 assign { out[138], out[394], out[650], out[906] } = in[111:108];
	 assign { out[137], out[393], out[649], out[905] } = in[119:116];
	 assign { out[136], out[392], out[648], out[904] } = in[127:124];
	 assign { out[151], out[407], out[663], out[919] } = in[135:132];
	 assign { out[150], out[406], out[662], out[918] } = in[143:140];
	 assign { out[149], out[405], out[661], out[917] } = in[151:148];
	 assign { out[148], out[404], out[660], out[916] } = in[159:156];
	 assign { out[147], out[403], out[659], out[915] } = in[167:164];
	 assign { out[146], out[402], out[658], out[914] } = in[175:172];
	 assign { out[145], out[401], out[657], out[913] } = in[183:180];
	 assign { out[144], out[400], out[656], out[912] } = in[191:188];
	 assign { out[159], out[415], out[671], out[927] } = in[199:196];
	 assign { out[158], out[414], out[670], out[926] } = in[207:204];
	 assign { out[157], out[413], out[669], out[925] } = in[215:212];
	 assign { out[156], out[412], out[668], out[924] } = in[223:220];
	 assign { out[155], out[411], out[667], out[923] } = in[231:228];
	 assign { out[154], out[410], out[666], out[922] } = in[239:236];
	 assign { out[153], out[409], out[665], out[921] } = in[247:244];
	 assign { out[152], out[408], out[664], out[920] } = in[255:252];
	 assign { out[167], out[423], out[679], out[935] } = in[263:260];
	 assign { out[166], out[422], out[678], out[934] } = in[271:268];
	 assign { out[165], out[421], out[677], out[933] } = in[279:276];
	 assign { out[164], out[420], out[676], out[932] } = in[287:284];
	 assign { out[163], out[419], out[675], out[931] } = in[295:292];
	 assign { out[162], out[418], out[674], out[930] } = in[303:300];
	 assign { out[161], out[417], out[673], out[929] } = in[311:308];
	 assign { out[160], out[416], out[672], out[928] } = in[319:316];
	 assign { out[175], out[431], out[687], out[943] } = in[327:324];
	 assign { out[174], out[430], out[686], out[942] } = in[335:332];
	 assign { out[173], out[429], out[685], out[941] } = in[343:340];
	 assign { out[172], out[428], out[684], out[940] } = in[351:348];
	 assign { out[171], out[427], out[683], out[939] } = in[359:356];
	 assign { out[170], out[426], out[682], out[938] } = in[367:364];
	 assign { out[169], out[425], out[681], out[937] } = in[375:372];
	 assign { out[168], out[424], out[680], out[936] } = in[383:380];
	 assign { out[183], out[439], out[695], out[951] } = in[391:388];
	 assign { out[182], out[438], out[694], out[950] } = in[399:396];
	 assign { out[181], out[437], out[693], out[949] } = in[407:404];
	 assign { out[180], out[436], out[692], out[948] } = in[415:412];
	 assign { out[179], out[435], out[691], out[947] } = in[423:420];
	 assign { out[178], out[434], out[690], out[946] } = in[431:428];
	 assign { out[177], out[433], out[689], out[945] } = in[439:436];
	 assign { out[176], out[432], out[688], out[944] } = in[447:444];
	 assign { out[191], out[447], out[703], out[959] } = in[455:452];
	 assign { out[190], out[446], out[702], out[958] } = in[463:460];
	 assign { out[189], out[445], out[701], out[957] } = in[471:468];
	 assign { out[188], out[444], out[700], out[956] } = in[479:476];
	 assign { out[187], out[443], out[699], out[955] } = in[487:484];
	 assign { out[186], out[442], out[698], out[954] } = in[495:492];
	 assign { out[185], out[441], out[697], out[953] } = in[503:500];
	 assign { out[184], out[440], out[696], out[952] } = in[511:508];
	 assign { out[199], out[455], out[711], out[967] } = in[519:516];
	 assign { out[198], out[454], out[710], out[966] } = in[527:524];
	 assign { out[197], out[453], out[709], out[965] } = in[535:532];
	 assign { out[196], out[452], out[708], out[964] } = in[543:540];
	 assign { out[195], out[451], out[707], out[963] } = in[551:548];
	 assign { out[194], out[450], out[706], out[962] } = in[559:556];
	 assign { out[193], out[449], out[705], out[961] } = in[567:564];
	 assign { out[192], out[448], out[704], out[960] } = in[575:572];
	 assign { out[207], out[463], out[719], out[975] } = in[583:580];
	 assign { out[206], out[462], out[718], out[974] } = in[591:588];
	 assign { out[205], out[461], out[717], out[973] } = in[599:596];
	 assign { out[204], out[460], out[716], out[972] } = in[607:604];
	 assign { out[203], out[459], out[715], out[971] } = in[615:612];
	 assign { out[202], out[458], out[714], out[970] } = in[623:620];
	 assign { out[201], out[457], out[713], out[969] } = in[631:628];
	 assign { out[200], out[456], out[712], out[968] } = in[639:636];
	 assign { out[215], out[471], out[727], out[983] } = in[647:644];
	 assign { out[214], out[470], out[726], out[982] } = in[655:652];
	 assign { out[213], out[469], out[725], out[981] } = in[663:660];
	 assign { out[212], out[468], out[724], out[980] } = in[671:668];
	 assign { out[211], out[467], out[723], out[979] } = in[679:676];
	 assign { out[210], out[466], out[722], out[978] } = in[687:684];
	 assign { out[209], out[465], out[721], out[977] } = in[695:692];
	 assign { out[208], out[464], out[720], out[976] } = in[703:700];
	 assign { out[223], out[479], out[735], out[991] } = in[711:708];
	 assign { out[222], out[478], out[734], out[990] } = in[719:716];
	 assign { out[221], out[477], out[733], out[989] } = in[727:724];
	 assign { out[220], out[476], out[732], out[988] } = in[735:732];
	 assign { out[219], out[475], out[731], out[987] } = in[743:740];
	 assign { out[218], out[474], out[730], out[986] } = in[751:748];
	 assign { out[217], out[473], out[729], out[985] } = in[759:756];
	 assign { out[216], out[472], out[728], out[984] } = in[767:764];
	 assign { out[231], out[487], out[743], out[999] } = in[775:772];
	 assign { out[230], out[486], out[742], out[998] } = in[783:780];
	 assign { out[229], out[485], out[741], out[997] } = in[791:788];
	 assign { out[228], out[484], out[740], out[996] } = in[799:796];
	 assign { out[227], out[483], out[739], out[995] } = in[807:804];
	 assign { out[226], out[482], out[738], out[994] } = in[815:812];
	 assign { out[225], out[481], out[737], out[993] } = in[823:820];
	 assign { out[224], out[480], out[736], out[992] } = in[831:828];
	 assign { out[239], out[495], out[751], out[1007] } = in[839:836];
	 assign { out[238], out[494], out[750], out[1006] } = in[847:844];
	 assign { out[237], out[493], out[749], out[1005] } = in[855:852];
	 assign { out[236], out[492], out[748], out[1004] } = in[863:860];
	 assign { out[235], out[491], out[747], out[1003] } = in[871:868];
	 assign { out[234], out[490], out[746], out[1002] } = in[879:876];
	 assign { out[233], out[489], out[745], out[1001] } = in[887:884];
	 assign { out[232], out[488], out[744], out[1000] } = in[895:892];
	 assign { out[247], out[503], out[759], out[1015] } = in[903:900];
	 assign { out[246], out[502], out[758], out[1014] } = in[911:908];
	 assign { out[245], out[501], out[757], out[1013] } = in[919:916];
	 assign { out[244], out[500], out[756], out[1012] } = in[927:924];
	 assign { out[243], out[499], out[755], out[1011] } = in[935:932];
	 assign { out[242], out[498], out[754], out[1010] } = in[943:940];
	 assign { out[241], out[497], out[753], out[1009] } = in[951:948];
	 assign { out[240], out[496], out[752], out[1008] } = in[959:956];
	 assign { out[255], out[511], out[767], out[1023] } = in[967:964];
	 assign { out[254], out[510], out[766], out[1022] } = in[975:972];
	 assign { out[253], out[509], out[765], out[1021] } = in[983:980];
	 assign { out[252], out[508], out[764], out[1020] } = in[991:988];
	 assign { out[251], out[507], out[763], out[1019] } = in[999:996];
	 assign { out[250], out[506], out[762], out[1018] } = in[1007:1004];
	 assign { out[249], out[505], out[761], out[1017] } = in[1015:1012];
	 assign { out[248], out[504], out[760], out[1016] } = in[1023:1020];

endmodule
